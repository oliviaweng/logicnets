module ens0_layer0 (input [783:0] M0, output [1023:0] M1);

wire [7:0] ens0_layer0_N0_wire = {M0[24], M0[72], M0[84], M0[315], M0[349], M0[435], M0[630], M0[724]};
ens0_layer0_N0 ens0_layer0_N0_inst (.M0(ens0_layer0_N0_wire), .M1(M1[0:0]));

wire [7:0] ens0_layer0_N1_wire = {M0[6], M0[267], M0[290], M0[362], M0[401], M0[434], M0[471], M0[579]};
ens0_layer0_N1 ens0_layer0_N1_inst (.M0(ens0_layer0_N1_wire), .M1(M1[1:1]));

wire [7:0] ens0_layer0_N2_wire = {M0[112], M0[117], M0[315], M0[332], M0[342], M0[366], M0[432], M0[606]};
ens0_layer0_N2 ens0_layer0_N2_inst (.M0(ens0_layer0_N2_wire), .M1(M1[2:2]));

wire [7:0] ens0_layer0_N3_wire = {M0[189], M0[277], M0[314], M0[400], M0[406], M0[576], M0[615], M0[625]};
ens0_layer0_N3 ens0_layer0_N3_inst (.M0(ens0_layer0_N3_wire), .M1(M1[3:3]));

wire [7:0] ens0_layer0_N4_wire = {M0[67], M0[132], M0[327], M0[441], M0[503], M0[716], M0[724], M0[759]};
ens0_layer0_N4 ens0_layer0_N4_inst (.M0(ens0_layer0_N4_wire), .M1(M1[4:4]));

wire [7:0] ens0_layer0_N5_wire = {M0[184], M0[285], M0[308], M0[311], M0[363], M0[442], M0[506], M0[545]};
ens0_layer0_N5 ens0_layer0_N5_inst (.M0(ens0_layer0_N5_wire), .M1(M1[5:5]));

wire [7:0] ens0_layer0_N6_wire = {M0[134], M0[330], M0[340], M0[448], M0[619], M0[640], M0[674], M0[686]};
ens0_layer0_N6 ens0_layer0_N6_inst (.M0(ens0_layer0_N6_wire), .M1(M1[6:6]));

wire [7:0] ens0_layer0_N7_wire = {M0[142], M0[186], M0[328], M0[341], M0[347], M0[395], M0[499], M0[662]};
ens0_layer0_N7 ens0_layer0_N7_inst (.M0(ens0_layer0_N7_wire), .M1(M1[7:7]));

wire [7:0] ens0_layer0_N8_wire = {M0[163], M0[172], M0[269], M0[349], M0[393], M0[424], M0[539], M0[689]};
ens0_layer0_N8 ens0_layer0_N8_inst (.M0(ens0_layer0_N8_wire), .M1(M1[8:8]));

wire [7:0] ens0_layer0_N9_wire = {M0[130], M0[309], M0[366], M0[410], M0[475], M0[518], M0[735], M0[762]};
ens0_layer0_N9 ens0_layer0_N9_inst (.M0(ens0_layer0_N9_wire), .M1(M1[9:9]));

wire [7:0] ens0_layer0_N10_wire = {M0[26], M0[58], M0[149], M0[429], M0[527], M0[559], M0[597], M0[621]};
ens0_layer0_N10 ens0_layer0_N10_inst (.M0(ens0_layer0_N10_wire), .M1(M1[10:10]));

wire [7:0] ens0_layer0_N11_wire = {M0[22], M0[84], M0[98], M0[203], M0[290], M0[312], M0[444], M0[691]};
ens0_layer0_N11 ens0_layer0_N11_inst (.M0(ens0_layer0_N11_wire), .M1(M1[11:11]));

wire [7:0] ens0_layer0_N12_wire = {M0[26], M0[65], M0[114], M0[369], M0[442], M0[525], M0[563], M0[622]};
ens0_layer0_N12 ens0_layer0_N12_inst (.M0(ens0_layer0_N12_wire), .M1(M1[12:12]));

wire [7:0] ens0_layer0_N13_wire = {M0[190], M0[251], M0[279], M0[401], M0[518], M0[621], M0[731], M0[760]};
ens0_layer0_N13 ens0_layer0_N13_inst (.M0(ens0_layer0_N13_wire), .M1(M1[13:13]));

wire [7:0] ens0_layer0_N14_wire = {M0[46], M0[132], M0[149], M0[249], M0[387], M0[507], M0[683], M0[750]};
ens0_layer0_N14 ens0_layer0_N14_inst (.M0(ens0_layer0_N14_wire), .M1(M1[14:14]));

wire [7:0] ens0_layer0_N15_wire = {M0[16], M0[148], M0[216], M0[310], M0[337], M0[364], M0[402], M0[634]};
ens0_layer0_N15 ens0_layer0_N15_inst (.M0(ens0_layer0_N15_wire), .M1(M1[15:15]));

wire [7:0] ens0_layer0_N16_wire = {M0[20], M0[76], M0[132], M0[185], M0[192], M0[345], M0[364], M0[466]};
ens0_layer0_N16 ens0_layer0_N16_inst (.M0(ens0_layer0_N16_wire), .M1(M1[16:16]));

wire [7:0] ens0_layer0_N17_wire = {M0[56], M0[97], M0[249], M0[358], M0[432], M0[433], M0[540], M0[551]};
ens0_layer0_N17 ens0_layer0_N17_inst (.M0(ens0_layer0_N17_wire), .M1(M1[17:17]));

wire [7:0] ens0_layer0_N18_wire = {M0[104], M0[174], M0[313], M0[425], M0[436], M0[621], M0[688], M0[729]};
ens0_layer0_N18 ens0_layer0_N18_inst (.M0(ens0_layer0_N18_wire), .M1(M1[18:18]));

wire [7:0] ens0_layer0_N19_wire = {M0[35], M0[230], M0[246], M0[360], M0[404], M0[525], M0[614], M0[748]};
ens0_layer0_N19 ens0_layer0_N19_inst (.M0(ens0_layer0_N19_wire), .M1(M1[19:19]));

wire [7:0] ens0_layer0_N20_wire = {M0[65], M0[364], M0[376], M0[483], M0[502], M0[507], M0[518], M0[661]};
ens0_layer0_N20 ens0_layer0_N20_inst (.M0(ens0_layer0_N20_wire), .M1(M1[20:20]));

wire [7:0] ens0_layer0_N21_wire = {M0[85], M0[242], M0[356], M0[542], M0[577], M0[702], M0[757], M0[776]};
ens0_layer0_N21 ens0_layer0_N21_inst (.M0(ens0_layer0_N21_wire), .M1(M1[21:21]));

wire [7:0] ens0_layer0_N22_wire = {M0[92], M0[254], M0[256], M0[267], M0[296], M0[531], M0[620], M0[663]};
ens0_layer0_N22 ens0_layer0_N22_inst (.M0(ens0_layer0_N22_wire), .M1(M1[22:22]));

wire [7:0] ens0_layer0_N23_wire = {M0[124], M0[215], M0[260], M0[362], M0[387], M0[436], M0[503], M0[617]};
ens0_layer0_N23 ens0_layer0_N23_inst (.M0(ens0_layer0_N23_wire), .M1(M1[23:23]));

wire [7:0] ens0_layer0_N24_wire = {M0[51], M0[97], M0[179], M0[195], M0[351], M0[360], M0[392], M0[622]};
ens0_layer0_N24 ens0_layer0_N24_inst (.M0(ens0_layer0_N24_wire), .M1(M1[24:24]));

wire [7:0] ens0_layer0_N25_wire = {M0[16], M0[293], M0[365], M0[406], M0[548], M0[575], M0[646], M0[783]};
ens0_layer0_N25 ens0_layer0_N25_inst (.M0(ens0_layer0_N25_wire), .M1(M1[25:25]));

wire [7:0] ens0_layer0_N26_wire = {M0[320], M0[391], M0[520], M0[524], M0[566], M0[654], M0[668], M0[687]};
ens0_layer0_N26 ens0_layer0_N26_inst (.M0(ens0_layer0_N26_wire), .M1(M1[26:26]));

wire [7:0] ens0_layer0_N27_wire = {M0[18], M0[46], M0[80], M0[86], M0[135], M0[277], M0[515], M0[529]};
ens0_layer0_N27 ens0_layer0_N27_inst (.M0(ens0_layer0_N27_wire), .M1(M1[27:27]));

wire [7:0] ens0_layer0_N28_wire = {M0[8], M0[111], M0[237], M0[266], M0[309], M0[384], M0[464], M0[754]};
ens0_layer0_N28 ens0_layer0_N28_inst (.M0(ens0_layer0_N28_wire), .M1(M1[28:28]));

wire [7:0] ens0_layer0_N29_wire = {M0[294], M0[396], M0[432], M0[483], M0[618], M0[635], M0[656], M0[701]};
ens0_layer0_N29 ens0_layer0_N29_inst (.M0(ens0_layer0_N29_wire), .M1(M1[29:29]));

wire [7:0] ens0_layer0_N30_wire = {M0[14], M0[66], M0[108], M0[379], M0[468], M0[586], M0[607], M0[649]};
ens0_layer0_N30 ens0_layer0_N30_inst (.M0(ens0_layer0_N30_wire), .M1(M1[30:30]));

wire [7:0] ens0_layer0_N31_wire = {M0[62], M0[170], M0[176], M0[197], M0[367], M0[383], M0[425], M0[655]};
ens0_layer0_N31 ens0_layer0_N31_inst (.M0(ens0_layer0_N31_wire), .M1(M1[31:31]));

wire [7:0] ens0_layer0_N32_wire = {M0[34], M0[342], M0[344], M0[369], M0[394], M0[613], M0[652], M0[656]};
ens0_layer0_N32 ens0_layer0_N32_inst (.M0(ens0_layer0_N32_wire), .M1(M1[32:32]));

wire [7:0] ens0_layer0_N33_wire = {M0[63], M0[398], M0[481], M0[493], M0[577], M0[692], M0[693], M0[719]};
ens0_layer0_N33 ens0_layer0_N33_inst (.M0(ens0_layer0_N33_wire), .M1(M1[33:33]));

wire [7:0] ens0_layer0_N34_wire = {M0[15], M0[78], M0[85], M0[174], M0[566], M0[622], M0[657], M0[774]};
ens0_layer0_N34 ens0_layer0_N34_inst (.M0(ens0_layer0_N34_wire), .M1(M1[34:34]));

wire [7:0] ens0_layer0_N35_wire = {M0[37], M0[84], M0[207], M0[222], M0[270], M0[279], M0[362], M0[389]};
ens0_layer0_N35 ens0_layer0_N35_inst (.M0(ens0_layer0_N35_wire), .M1(M1[35:35]));

wire [7:0] ens0_layer0_N36_wire = {M0[47], M0[165], M0[333], M0[375], M0[411], M0[424], M0[624], M0[777]};
ens0_layer0_N36 ens0_layer0_N36_inst (.M0(ens0_layer0_N36_wire), .M1(M1[36:36]));

wire [7:0] ens0_layer0_N37_wire = {M0[56], M0[172], M0[231], M0[382], M0[432], M0[533], M0[536], M0[647]};
ens0_layer0_N37 ens0_layer0_N37_inst (.M0(ens0_layer0_N37_wire), .M1(M1[37:37]));

wire [7:0] ens0_layer0_N38_wire = {M0[66], M0[132], M0[215], M0[307], M0[328], M0[408], M0[680], M0[740]};
ens0_layer0_N38 ens0_layer0_N38_inst (.M0(ens0_layer0_N38_wire), .M1(M1[38:38]));

wire [7:0] ens0_layer0_N39_wire = {M0[285], M0[290], M0[435], M0[451], M0[475], M0[539], M0[606], M0[624]};
ens0_layer0_N39 ens0_layer0_N39_inst (.M0(ens0_layer0_N39_wire), .M1(M1[39:39]));

wire [7:0] ens0_layer0_N40_wire = {M0[46], M0[132], M0[169], M0[393], M0[442], M0[616], M0[702], M0[772]};
ens0_layer0_N40 ens0_layer0_N40_inst (.M0(ens0_layer0_N40_wire), .M1(M1[40:40]));

wire [7:0] ens0_layer0_N41_wire = {M0[152], M0[207], M0[360], M0[420], M0[514], M0[544], M0[548], M0[667]};
ens0_layer0_N41 ens0_layer0_N41_inst (.M0(ens0_layer0_N41_wire), .M1(M1[41:41]));

wire [7:0] ens0_layer0_N42_wire = {M0[103], M0[268], M0[306], M0[342], M0[497], M0[501], M0[548], M0[684]};
ens0_layer0_N42 ens0_layer0_N42_inst (.M0(ens0_layer0_N42_wire), .M1(M1[42:42]));

wire [7:0] ens0_layer0_N43_wire = {M0[142], M0[320], M0[363], M0[378], M0[523], M0[525], M0[749], M0[776]};
ens0_layer0_N43 ens0_layer0_N43_inst (.M0(ens0_layer0_N43_wire), .M1(M1[43:43]));

wire [7:0] ens0_layer0_N44_wire = {M0[288], M0[331], M0[457], M0[468], M0[648], M0[664], M0[678], M0[760]};
ens0_layer0_N44 ens0_layer0_N44_inst (.M0(ens0_layer0_N44_wire), .M1(M1[44:44]));

wire [7:0] ens0_layer0_N45_wire = {M0[13], M0[178], M0[413], M0[450], M0[467], M0[512], M0[660], M0[777]};
ens0_layer0_N45 ens0_layer0_N45_inst (.M0(ens0_layer0_N45_wire), .M1(M1[45:45]));

wire [7:0] ens0_layer0_N46_wire = {M0[178], M0[225], M0[306], M0[350], M0[441], M0[612], M0[649], M0[671]};
ens0_layer0_N46 ens0_layer0_N46_inst (.M0(ens0_layer0_N46_wire), .M1(M1[46:46]));

wire [7:0] ens0_layer0_N47_wire = {M0[164], M0[201], M0[270], M0[530], M0[554], M0[555], M0[612], M0[725]};
ens0_layer0_N47 ens0_layer0_N47_inst (.M0(ens0_layer0_N47_wire), .M1(M1[47:47]));

wire [7:0] ens0_layer0_N48_wire = {M0[17], M0[184], M0[212], M0[331], M0[470], M0[533], M0[694], M0[717]};
ens0_layer0_N48 ens0_layer0_N48_inst (.M0(ens0_layer0_N48_wire), .M1(M1[48:48]));

wire [7:0] ens0_layer0_N49_wire = {M0[62], M0[79], M0[172], M0[339], M0[423], M0[556], M0[649], M0[721]};
ens0_layer0_N49 ens0_layer0_N49_inst (.M0(ens0_layer0_N49_wire), .M1(M1[49:49]));

wire [7:0] ens0_layer0_N50_wire = {M0[65], M0[321], M0[371], M0[387], M0[537], M0[582], M0[641], M0[661]};
ens0_layer0_N50 ens0_layer0_N50_inst (.M0(ens0_layer0_N50_wire), .M1(M1[50:50]));

wire [7:0] ens0_layer0_N51_wire = {M0[297], M0[355], M0[496], M0[535], M0[556], M0[649], M0[653], M0[713]};
ens0_layer0_N51 ens0_layer0_N51_inst (.M0(ens0_layer0_N51_wire), .M1(M1[51:51]));

wire [7:0] ens0_layer0_N52_wire = {M0[71], M0[205], M0[391], M0[615], M0[629], M0[679], M0[703], M0[772]};
ens0_layer0_N52 ens0_layer0_N52_inst (.M0(ens0_layer0_N52_wire), .M1(M1[52:52]));

wire [7:0] ens0_layer0_N53_wire = {M0[48], M0[113], M0[116], M0[389], M0[502], M0[655], M0[713], M0[714]};
ens0_layer0_N53 ens0_layer0_N53_inst (.M0(ens0_layer0_N53_wire), .M1(M1[53:53]));

wire [7:0] ens0_layer0_N54_wire = {M0[154], M0[172], M0[282], M0[392], M0[541], M0[570], M0[642], M0[781]};
ens0_layer0_N54 ens0_layer0_N54_inst (.M0(ens0_layer0_N54_wire), .M1(M1[54:54]));

wire [7:0] ens0_layer0_N55_wire = {M0[163], M0[191], M0[246], M0[317], M0[356], M0[495], M0[511], M0[548]};
ens0_layer0_N55 ens0_layer0_N55_inst (.M0(ens0_layer0_N55_wire), .M1(M1[55:55]));

wire [7:0] ens0_layer0_N56_wire = {M0[41], M0[52], M0[59], M0[129], M0[146], M0[260], M0[565], M0[682]};
ens0_layer0_N56 ens0_layer0_N56_inst (.M0(ens0_layer0_N56_wire), .M1(M1[56:56]));

wire [7:0] ens0_layer0_N57_wire = {M0[27], M0[184], M0[216], M0[244], M0[247], M0[414], M0[658], M0[783]};
ens0_layer0_N57 ens0_layer0_N57_inst (.M0(ens0_layer0_N57_wire), .M1(M1[57:57]));

wire [7:0] ens0_layer0_N58_wire = {M0[179], M0[195], M0[366], M0[506], M0[625], M0[683], M0[743], M0[780]};
ens0_layer0_N58 ens0_layer0_N58_inst (.M0(ens0_layer0_N58_wire), .M1(M1[58:58]));

wire [7:0] ens0_layer0_N59_wire = {M0[156], M0[239], M0[263], M0[338], M0[359], M0[723], M0[724], M0[729]};
ens0_layer0_N59 ens0_layer0_N59_inst (.M0(ens0_layer0_N59_wire), .M1(M1[59:59]));

wire [7:0] ens0_layer0_N60_wire = {M0[11], M0[108], M0[113], M0[334], M0[391], M0[538], M0[639], M0[764]};
ens0_layer0_N60 ens0_layer0_N60_inst (.M0(ens0_layer0_N60_wire), .M1(M1[60:60]));

wire [7:0] ens0_layer0_N61_wire = {M0[42], M0[292], M0[314], M0[363], M0[636], M0[663], M0[671], M0[755]};
ens0_layer0_N61 ens0_layer0_N61_inst (.M0(ens0_layer0_N61_wire), .M1(M1[61:61]));

wire [7:0] ens0_layer0_N62_wire = {M0[35], M0[64], M0[221], M0[228], M0[487], M0[562], M0[564], M0[623]};
ens0_layer0_N62 ens0_layer0_N62_inst (.M0(ens0_layer0_N62_wire), .M1(M1[62:62]));

wire [7:0] ens0_layer0_N63_wire = {M0[93], M0[145], M0[236], M0[246], M0[456], M0[740], M0[744], M0[766]};
ens0_layer0_N63 ens0_layer0_N63_inst (.M0(ens0_layer0_N63_wire), .M1(M1[63:63]));

wire [7:0] ens0_layer0_N64_wire = {M0[3], M0[342], M0[387], M0[409], M0[431], M0[610], M0[683], M0[737]};
ens0_layer0_N64 ens0_layer0_N64_inst (.M0(ens0_layer0_N64_wire), .M1(M1[64:64]));

wire [7:0] ens0_layer0_N65_wire = {M0[60], M0[124], M0[195], M0[207], M0[223], M0[255], M0[410], M0[567]};
ens0_layer0_N65 ens0_layer0_N65_inst (.M0(ens0_layer0_N65_wire), .M1(M1[65:65]));

wire [7:0] ens0_layer0_N66_wire = {M0[11], M0[89], M0[97], M0[234], M0[509], M0[526], M0[633], M0[645]};
ens0_layer0_N66 ens0_layer0_N66_inst (.M0(ens0_layer0_N66_wire), .M1(M1[66:66]));

wire [7:0] ens0_layer0_N67_wire = {M0[44], M0[195], M0[243], M0[349], M0[450], M0[480], M0[551], M0[651]};
ens0_layer0_N67 ens0_layer0_N67_inst (.M0(ens0_layer0_N67_wire), .M1(M1[67:67]));

wire [7:0] ens0_layer0_N68_wire = {M0[8], M0[9], M0[271], M0[304], M0[554], M0[651], M0[663], M0[782]};
ens0_layer0_N68 ens0_layer0_N68_inst (.M0(ens0_layer0_N68_wire), .M1(M1[68:68]));

wire [7:0] ens0_layer0_N69_wire = {M0[27], M0[166], M0[174], M0[180], M0[199], M0[304], M0[629], M0[707]};
ens0_layer0_N69 ens0_layer0_N69_inst (.M0(ens0_layer0_N69_wire), .M1(M1[69:69]));

wire [7:0] ens0_layer0_N70_wire = {M0[3], M0[17], M0[261], M0[439], M0[528], M0[648], M0[664], M0[770]};
ens0_layer0_N70 ens0_layer0_N70_inst (.M0(ens0_layer0_N70_wire), .M1(M1[70:70]));

wire [7:0] ens0_layer0_N71_wire = {M0[27], M0[118], M0[267], M0[446], M0[511], M0[557], M0[561], M0[580]};
ens0_layer0_N71 ens0_layer0_N71_inst (.M0(ens0_layer0_N71_wire), .M1(M1[71:71]));

wire [7:0] ens0_layer0_N72_wire = {M0[43], M0[234], M0[377], M0[448], M0[663], M0[689], M0[715], M0[749]};
ens0_layer0_N72 ens0_layer0_N72_inst (.M0(ens0_layer0_N72_wire), .M1(M1[72:72]));

wire [7:0] ens0_layer0_N73_wire = {M0[56], M0[261], M0[350], M0[450], M0[482], M0[566], M0[654], M0[692]};
ens0_layer0_N73 ens0_layer0_N73_inst (.M0(ens0_layer0_N73_wire), .M1(M1[73:73]));

wire [7:0] ens0_layer0_N74_wire = {M0[166], M0[205], M0[479], M0[496], M0[531], M0[552], M0[618], M0[677]};
ens0_layer0_N74 ens0_layer0_N74_inst (.M0(ens0_layer0_N74_wire), .M1(M1[74:74]));

wire [7:0] ens0_layer0_N75_wire = {M0[10], M0[266], M0[390], M0[396], M0[397], M0[459], M0[649], M0[773]};
ens0_layer0_N75 ens0_layer0_N75_inst (.M0(ens0_layer0_N75_wire), .M1(M1[75:75]));

wire [7:0] ens0_layer0_N76_wire = {M0[54], M0[252], M0[340], M0[359], M0[473], M0[524], M0[666], M0[757]};
ens0_layer0_N76 ens0_layer0_N76_inst (.M0(ens0_layer0_N76_wire), .M1(M1[76:76]));

wire [7:0] ens0_layer0_N77_wire = {M0[0], M0[114], M0[190], M0[253], M0[257], M0[442], M0[504], M0[702]};
ens0_layer0_N77 ens0_layer0_N77_inst (.M0(ens0_layer0_N77_wire), .M1(M1[77:77]));

wire [7:0] ens0_layer0_N78_wire = {M0[154], M0[298], M0[326], M0[328], M0[435], M0[593], M0[686], M0[709]};
ens0_layer0_N78 ens0_layer0_N78_inst (.M0(ens0_layer0_N78_wire), .M1(M1[78:78]));

wire [7:0] ens0_layer0_N79_wire = {M0[171], M0[293], M0[300], M0[406], M0[552], M0[605], M0[655], M0[764]};
ens0_layer0_N79 ens0_layer0_N79_inst (.M0(ens0_layer0_N79_wire), .M1(M1[79:79]));

wire [7:0] ens0_layer0_N80_wire = {M0[96], M0[150], M0[178], M0[252], M0[369], M0[615], M0[686], M0[783]};
ens0_layer0_N80 ens0_layer0_N80_inst (.M0(ens0_layer0_N80_wire), .M1(M1[80:80]));

wire [7:0] ens0_layer0_N81_wire = {M0[10], M0[101], M0[189], M0[449], M0[525], M0[564], M0[626], M0[642]};
ens0_layer0_N81 ens0_layer0_N81_inst (.M0(ens0_layer0_N81_wire), .M1(M1[81:81]));

wire [7:0] ens0_layer0_N82_wire = {M0[21], M0[34], M0[133], M0[177], M0[180], M0[620], M0[657], M0[776]};
ens0_layer0_N82 ens0_layer0_N82_inst (.M0(ens0_layer0_N82_wire), .M1(M1[82:82]));

wire [7:0] ens0_layer0_N83_wire = {M0[13], M0[310], M0[499], M0[531], M0[540], M0[640], M0[691], M0[702]};
ens0_layer0_N83 ens0_layer0_N83_inst (.M0(ens0_layer0_N83_wire), .M1(M1[83:83]));

wire [7:0] ens0_layer0_N84_wire = {M0[92], M0[279], M0[287], M0[466], M0[484], M0[520], M0[577], M0[622]};
ens0_layer0_N84 ens0_layer0_N84_inst (.M0(ens0_layer0_N84_wire), .M1(M1[84:84]));

wire [7:0] ens0_layer0_N85_wire = {M0[64], M0[175], M0[256], M0[358], M0[413], M0[434], M0[638], M0[679]};
ens0_layer0_N85 ens0_layer0_N85_inst (.M0(ens0_layer0_N85_wire), .M1(M1[85:85]));

wire [7:0] ens0_layer0_N86_wire = {M0[116], M0[131], M0[199], M0[367], M0[617], M0[652], M0[731], M0[741]};
ens0_layer0_N86 ens0_layer0_N86_inst (.M0(ens0_layer0_N86_wire), .M1(M1[86:86]));

wire [7:0] ens0_layer0_N87_wire = {M0[68], M0[208], M0[213], M0[429], M0[462], M0[495], M0[544], M0[767]};
ens0_layer0_N87 ens0_layer0_N87_inst (.M0(ens0_layer0_N87_wire), .M1(M1[87:87]));

wire [7:0] ens0_layer0_N88_wire = {M0[127], M0[278], M0[414], M0[526], M0[531], M0[548], M0[637], M0[658]};
ens0_layer0_N88 ens0_layer0_N88_inst (.M0(ens0_layer0_N88_wire), .M1(M1[88:88]));

wire [7:0] ens0_layer0_N89_wire = {M0[327], M0[328], M0[439], M0[525], M0[562], M0[566], M0[606], M0[668]};
ens0_layer0_N89 ens0_layer0_N89_inst (.M0(ens0_layer0_N89_wire), .M1(M1[89:89]));

wire [7:0] ens0_layer0_N90_wire = {M0[9], M0[224], M0[234], M0[294], M0[387], M0[512], M0[541], M0[588]};
ens0_layer0_N90 ens0_layer0_N90_inst (.M0(ens0_layer0_N90_wire), .M1(M1[90:90]));

wire [7:0] ens0_layer0_N91_wire = {M0[56], M0[197], M0[600], M0[604], M0[697], M0[700], M0[719], M0[768]};
ens0_layer0_N91 ens0_layer0_N91_inst (.M0(ens0_layer0_N91_wire), .M1(M1[91:91]));

wire [7:0] ens0_layer0_N92_wire = {M0[188], M0[226], M0[245], M0[400], M0[497], M0[628], M0[677], M0[778]};
ens0_layer0_N92 ens0_layer0_N92_inst (.M0(ens0_layer0_N92_wire), .M1(M1[92:92]));

wire [7:0] ens0_layer0_N93_wire = {M0[69], M0[185], M0[402], M0[424], M0[473], M0[474], M0[560], M0[640]};
ens0_layer0_N93 ens0_layer0_N93_inst (.M0(ens0_layer0_N93_wire), .M1(M1[93:93]));

wire [7:0] ens0_layer0_N94_wire = {M0[21], M0[38], M0[111], M0[140], M0[163], M0[244], M0[443], M0[486]};
ens0_layer0_N94 ens0_layer0_N94_inst (.M0(ens0_layer0_N94_wire), .M1(M1[94:94]));

wire [7:0] ens0_layer0_N95_wire = {M0[201], M0[206], M0[263], M0[378], M0[379], M0[426], M0[534], M0[644]};
ens0_layer0_N95 ens0_layer0_N95_inst (.M0(ens0_layer0_N95_wire), .M1(M1[95:95]));

wire [7:0] ens0_layer0_N96_wire = {M0[55], M0[132], M0[146], M0[261], M0[280], M0[489], M0[643], M0[765]};
ens0_layer0_N96 ens0_layer0_N96_inst (.M0(ens0_layer0_N96_wire), .M1(M1[96:96]));

wire [7:0] ens0_layer0_N97_wire = {M0[48], M0[71], M0[84], M0[299], M0[532], M0[561], M0[577], M0[708]};
ens0_layer0_N97 ens0_layer0_N97_inst (.M0(ens0_layer0_N97_wire), .M1(M1[97:97]));

wire [7:0] ens0_layer0_N98_wire = {M0[113], M0[304], M0[347], M0[384], M0[492], M0[560], M0[741], M0[772]};
ens0_layer0_N98 ens0_layer0_N98_inst (.M0(ens0_layer0_N98_wire), .M1(M1[98:98]));

wire [7:0] ens0_layer0_N99_wire = {M0[132], M0[260], M0[452], M0[467], M0[542], M0[733], M0[772], M0[779]};
ens0_layer0_N99 ens0_layer0_N99_inst (.M0(ens0_layer0_N99_wire), .M1(M1[99:99]));

wire [7:0] ens0_layer0_N100_wire = {M0[85], M0[258], M0[351], M0[444], M0[464], M0[500], M0[701], M0[752]};
ens0_layer0_N100 ens0_layer0_N100_inst (.M0(ens0_layer0_N100_wire), .M1(M1[100:100]));

wire [7:0] ens0_layer0_N101_wire = {M0[81], M0[95], M0[110], M0[245], M0[420], M0[651], M0[704], M0[783]};
ens0_layer0_N101 ens0_layer0_N101_inst (.M0(ens0_layer0_N101_wire), .M1(M1[101:101]));

wire [7:0] ens0_layer0_N102_wire = {M0[53], M0[84], M0[98], M0[351], M0[420], M0[528], M0[565], M0[723]};
ens0_layer0_N102 ens0_layer0_N102_inst (.M0(ens0_layer0_N102_wire), .M1(M1[102:102]));

wire [7:0] ens0_layer0_N103_wire = {M0[66], M0[171], M0[195], M0[290], M0[525], M0[647], M0[739], M0[780]};
ens0_layer0_N103 ens0_layer0_N103_inst (.M0(ens0_layer0_N103_wire), .M1(M1[103:103]));

wire [7:0] ens0_layer0_N104_wire = {M0[6], M0[64], M0[88], M0[292], M0[314], M0[398], M0[427], M0[565]};
ens0_layer0_N104 ens0_layer0_N104_inst (.M0(ens0_layer0_N104_wire), .M1(M1[104:104]));

wire [7:0] ens0_layer0_N105_wire = {M0[65], M0[127], M0[138], M0[193], M0[268], M0[274], M0[387], M0[645]};
ens0_layer0_N105 ens0_layer0_N105_inst (.M0(ens0_layer0_N105_wire), .M1(M1[105:105]));

wire [7:0] ens0_layer0_N106_wire = {M0[5], M0[78], M0[263], M0[345], M0[356], M0[402], M0[503], M0[554]};
ens0_layer0_N106 ens0_layer0_N106_inst (.M0(ens0_layer0_N106_wire), .M1(M1[106:106]));

wire [7:0] ens0_layer0_N107_wire = {M0[49], M0[66], M0[144], M0[177], M0[391], M0[412], M0[502], M0[625]};
ens0_layer0_N107 ens0_layer0_N107_inst (.M0(ens0_layer0_N107_wire), .M1(M1[107:107]));

wire [7:0] ens0_layer0_N108_wire = {M0[33], M0[286], M0[293], M0[424], M0[484], M0[517], M0[532], M0[739]};
ens0_layer0_N108 ens0_layer0_N108_inst (.M0(ens0_layer0_N108_wire), .M1(M1[108:108]));

wire [7:0] ens0_layer0_N109_wire = {M0[205], M0[249], M0[318], M0[327], M0[340], M0[387], M0[524], M0[672]};
ens0_layer0_N109 ens0_layer0_N109_inst (.M0(ens0_layer0_N109_wire), .M1(M1[109:109]));

wire [7:0] ens0_layer0_N110_wire = {M0[177], M0[222], M0[273], M0[291], M0[551], M0[557], M0[695], M0[768]};
ens0_layer0_N110 ens0_layer0_N110_inst (.M0(ens0_layer0_N110_wire), .M1(M1[110:110]));

wire [7:0] ens0_layer0_N111_wire = {M0[209], M0[285], M0[308], M0[461], M0[534], M0[554], M0[572], M0[717]};
ens0_layer0_N111 ens0_layer0_N111_inst (.M0(ens0_layer0_N111_wire), .M1(M1[111:111]));

wire [7:0] ens0_layer0_N112_wire = {M0[235], M0[239], M0[347], M0[437], M0[443], M0[446], M0[469], M0[610]};
ens0_layer0_N112 ens0_layer0_N112_inst (.M0(ens0_layer0_N112_wire), .M1(M1[112:112]));

wire [7:0] ens0_layer0_N113_wire = {M0[113], M0[247], M0[248], M0[325], M0[461], M0[466], M0[612], M0[759]};
ens0_layer0_N113 ens0_layer0_N113_inst (.M0(ens0_layer0_N113_wire), .M1(M1[113:113]));

wire [7:0] ens0_layer0_N114_wire = {M0[117], M0[205], M0[318], M0[560], M0[607], M0[617], M0[651], M0[722]};
ens0_layer0_N114 ens0_layer0_N114_inst (.M0(ens0_layer0_N114_wire), .M1(M1[114:114]));

wire [7:0] ens0_layer0_N115_wire = {M0[158], M0[169], M0[197], M0[308], M0[414], M0[463], M0[509], M0[512]};
ens0_layer0_N115 ens0_layer0_N115_inst (.M0(ens0_layer0_N115_wire), .M1(M1[115:115]));

wire [7:0] ens0_layer0_N116_wire = {M0[250], M0[404], M0[431], M0[441], M0[503], M0[660], M0[756], M0[768]};
ens0_layer0_N116 ens0_layer0_N116_inst (.M0(ens0_layer0_N116_wire), .M1(M1[116:116]));

wire [7:0] ens0_layer0_N117_wire = {M0[14], M0[133], M0[162], M0[310], M0[422], M0[528], M0[595], M0[738]};
ens0_layer0_N117 ens0_layer0_N117_inst (.M0(ens0_layer0_N117_wire), .M1(M1[117:117]));

wire [7:0] ens0_layer0_N118_wire = {M0[41], M0[90], M0[458], M0[533], M0[566], M0[567], M0[666], M0[711]};
ens0_layer0_N118 ens0_layer0_N118_inst (.M0(ens0_layer0_N118_wire), .M1(M1[118:118]));

wire [7:0] ens0_layer0_N119_wire = {M0[9], M0[44], M0[175], M0[180], M0[219], M0[322], M0[537], M0[757]};
ens0_layer0_N119 ens0_layer0_N119_inst (.M0(ens0_layer0_N119_wire), .M1(M1[119:119]));

wire [7:0] ens0_layer0_N120_wire = {M0[73], M0[153], M0[321], M0[332], M0[528], M0[533], M0[561], M0[745]};
ens0_layer0_N120 ens0_layer0_N120_inst (.M0(ens0_layer0_N120_wire), .M1(M1[120:120]));

wire [7:0] ens0_layer0_N121_wire = {M0[15], M0[46], M0[73], M0[117], M0[350], M0[688], M0[738], M0[751]};
ens0_layer0_N121 ens0_layer0_N121_inst (.M0(ens0_layer0_N121_wire), .M1(M1[121:121]));

wire [7:0] ens0_layer0_N122_wire = {M0[2], M0[60], M0[345], M0[435], M0[453], M0[741], M0[745], M0[778]};
ens0_layer0_N122 ens0_layer0_N122_inst (.M0(ens0_layer0_N122_wire), .M1(M1[122:122]));

wire [7:0] ens0_layer0_N123_wire = {M0[39], M0[156], M0[338], M0[456], M0[495], M0[508], M0[530], M0[728]};
ens0_layer0_N123 ens0_layer0_N123_inst (.M0(ens0_layer0_N123_wire), .M1(M1[123:123]));

wire [7:0] ens0_layer0_N124_wire = {M0[25], M0[109], M0[138], M0[181], M0[355], M0[393], M0[705], M0[718]};
ens0_layer0_N124 ens0_layer0_N124_inst (.M0(ens0_layer0_N124_wire), .M1(M1[124:124]));

wire [7:0] ens0_layer0_N125_wire = {M0[212], M0[290], M0[338], M0[378], M0[451], M0[474], M0[494], M0[634]};
ens0_layer0_N125 ens0_layer0_N125_inst (.M0(ens0_layer0_N125_wire), .M1(M1[125:125]));

wire [7:0] ens0_layer0_N126_wire = {M0[155], M0[227], M0[325], M0[457], M0[486], M0[535], M0[729], M0[732]};
ens0_layer0_N126 ens0_layer0_N126_inst (.M0(ens0_layer0_N126_wire), .M1(M1[126:126]));

wire [7:0] ens0_layer0_N127_wire = {M0[134], M0[180], M0[225], M0[257], M0[463], M0[606], M0[621], M0[757]};
ens0_layer0_N127 ens0_layer0_N127_inst (.M0(ens0_layer0_N127_wire), .M1(M1[127:127]));

wire [7:0] ens0_layer0_N128_wire = {M0[36], M0[349], M0[418], M0[487], M0[550], M0[558], M0[578], M0[731]};
ens0_layer0_N128 ens0_layer0_N128_inst (.M0(ens0_layer0_N128_wire), .M1(M1[128:128]));

wire [7:0] ens0_layer0_N129_wire = {M0[4], M0[57], M0[72], M0[209], M0[314], M0[490], M0[697], M0[733]};
ens0_layer0_N129 ens0_layer0_N129_inst (.M0(ens0_layer0_N129_wire), .M1(M1[129:129]));

wire [7:0] ens0_layer0_N130_wire = {M0[152], M0[217], M0[241], M0[274], M0[286], M0[328], M0[502], M0[777]};
ens0_layer0_N130 ens0_layer0_N130_inst (.M0(ens0_layer0_N130_wire), .M1(M1[130:130]));

wire [7:0] ens0_layer0_N131_wire = {M0[85], M0[112], M0[148], M0[281], M0[283], M0[311], M0[576], M0[724]};
ens0_layer0_N131 ens0_layer0_N131_inst (.M0(ens0_layer0_N131_wire), .M1(M1[131:131]));

wire [7:0] ens0_layer0_N132_wire = {M0[18], M0[43], M0[55], M0[111], M0[150], M0[260], M0[261], M0[489]};
ens0_layer0_N132 ens0_layer0_N132_inst (.M0(ens0_layer0_N132_wire), .M1(M1[132:132]));

wire [7:0] ens0_layer0_N133_wire = {M0[93], M0[290], M0[367], M0[422], M0[455], M0[573], M0[637], M0[641]};
ens0_layer0_N133 ens0_layer0_N133_inst (.M0(ens0_layer0_N133_wire), .M1(M1[133:133]));

wire [7:0] ens0_layer0_N134_wire = {M0[156], M0[193], M0[287], M0[332], M0[526], M0[551], M0[639], M0[683]};
ens0_layer0_N134 ens0_layer0_N134_inst (.M0(ens0_layer0_N134_wire), .M1(M1[134:134]));

wire [7:0] ens0_layer0_N135_wire = {M0[61], M0[129], M0[265], M0[326], M0[372], M0[378], M0[558], M0[666]};
ens0_layer0_N135 ens0_layer0_N135_inst (.M0(ens0_layer0_N135_wire), .M1(M1[135:135]));

wire [7:0] ens0_layer0_N136_wire = {M0[58], M0[291], M0[407], M0[448], M0[567], M0[629], M0[733], M0[774]};
ens0_layer0_N136 ens0_layer0_N136_inst (.M0(ens0_layer0_N136_wire), .M1(M1[136:136]));

wire [7:0] ens0_layer0_N137_wire = {M0[74], M0[172], M0[262], M0[269], M0[309], M0[477], M0[685], M0[745]};
ens0_layer0_N137 ens0_layer0_N137_inst (.M0(ens0_layer0_N137_wire), .M1(M1[137:137]));

wire [7:0] ens0_layer0_N138_wire = {M0[48], M0[115], M0[257], M0[294], M0[521], M0[612], M0[655], M0[770]};
ens0_layer0_N138 ens0_layer0_N138_inst (.M0(ens0_layer0_N138_wire), .M1(M1[138:138]));

wire [7:0] ens0_layer0_N139_wire = {M0[154], M0[191], M0[299], M0[349], M0[479], M0[586], M0[643], M0[683]};
ens0_layer0_N139 ens0_layer0_N139_inst (.M0(ens0_layer0_N139_wire), .M1(M1[139:139]));

wire [7:0] ens0_layer0_N140_wire = {M0[110], M0[273], M0[418], M0[454], M0[547], M0[551], M0[763], M0[780]};
ens0_layer0_N140 ens0_layer0_N140_inst (.M0(ens0_layer0_N140_wire), .M1(M1[140:140]));

wire [7:0] ens0_layer0_N141_wire = {M0[78], M0[154], M0[205], M0[406], M0[454], M0[579], M0[737], M0[770]};
ens0_layer0_N141 ens0_layer0_N141_inst (.M0(ens0_layer0_N141_wire), .M1(M1[141:141]));

wire [7:0] ens0_layer0_N142_wire = {M0[86], M0[339], M0[408], M0[409], M0[498], M0[521], M0[575], M0[645]};
ens0_layer0_N142 ens0_layer0_N142_inst (.M0(ens0_layer0_N142_wire), .M1(M1[142:142]));

wire [7:0] ens0_layer0_N143_wire = {M0[85], M0[237], M0[270], M0[305], M0[357], M0[452], M0[566], M0[718]};
ens0_layer0_N143 ens0_layer0_N143_inst (.M0(ens0_layer0_N143_wire), .M1(M1[143:143]));

wire [7:0] ens0_layer0_N144_wire = {M0[99], M0[200], M0[321], M0[391], M0[519], M0[666], M0[681], M0[692]};
ens0_layer0_N144 ens0_layer0_N144_inst (.M0(ens0_layer0_N144_wire), .M1(M1[144:144]));

wire [7:0] ens0_layer0_N145_wire = {M0[126], M0[160], M0[248], M0[324], M0[326], M0[442], M0[451], M0[763]};
ens0_layer0_N145 ens0_layer0_N145_inst (.M0(ens0_layer0_N145_wire), .M1(M1[145:145]));

wire [7:0] ens0_layer0_N146_wire = {M0[106], M0[134], M0[320], M0[474], M0[486], M0[518], M0[576], M0[628]};
ens0_layer0_N146 ens0_layer0_N146_inst (.M0(ens0_layer0_N146_wire), .M1(M1[146:146]));

wire [7:0] ens0_layer0_N147_wire = {M0[6], M0[135], M0[179], M0[214], M0[255], M0[348], M0[350], M0[490]};
ens0_layer0_N147 ens0_layer0_N147_inst (.M0(ens0_layer0_N147_wire), .M1(M1[147:147]));

wire [7:0] ens0_layer0_N148_wire = {M0[32], M0[133], M0[188], M0[226], M0[388], M0[442], M0[535], M0[690]};
ens0_layer0_N148 ens0_layer0_N148_inst (.M0(ens0_layer0_N148_wire), .M1(M1[148:148]));

wire [7:0] ens0_layer0_N149_wire = {M0[11], M0[105], M0[352], M0[412], M0[455], M0[565], M0[578], M0[649]};
ens0_layer0_N149 ens0_layer0_N149_inst (.M0(ens0_layer0_N149_wire), .M1(M1[149:149]));

wire [7:0] ens0_layer0_N150_wire = {M0[95], M0[136], M0[141], M0[174], M0[191], M0[491], M0[513], M0[616]};
ens0_layer0_N150 ens0_layer0_N150_inst (.M0(ens0_layer0_N150_wire), .M1(M1[150:150]));

wire [7:0] ens0_layer0_N151_wire = {M0[33], M0[294], M0[380], M0[582], M0[584], M0[621], M0[666], M0[771]};
ens0_layer0_N151 ens0_layer0_N151_inst (.M0(ens0_layer0_N151_wire), .M1(M1[151:151]));

wire [7:0] ens0_layer0_N152_wire = {M0[25], M0[71], M0[292], M0[380], M0[426], M0[475], M0[632], M0[664]};
ens0_layer0_N152 ens0_layer0_N152_inst (.M0(ens0_layer0_N152_wire), .M1(M1[152:152]));

wire [7:0] ens0_layer0_N153_wire = {M0[115], M0[238], M0[254], M0[294], M0[324], M0[359], M0[411], M0[750]};
ens0_layer0_N153 ens0_layer0_N153_inst (.M0(ens0_layer0_N153_wire), .M1(M1[153:153]));

wire [7:0] ens0_layer0_N154_wire = {M0[8], M0[72], M0[207], M0[275], M0[495], M0[587], M0[591], M0[745]};
ens0_layer0_N154 ens0_layer0_N154_inst (.M0(ens0_layer0_N154_wire), .M1(M1[154:154]));

wire [7:0] ens0_layer0_N155_wire = {M0[20], M0[270], M0[366], M0[396], M0[407], M0[500], M0[548], M0[717]};
ens0_layer0_N155 ens0_layer0_N155_inst (.M0(ens0_layer0_N155_wire), .M1(M1[155:155]));

wire [7:0] ens0_layer0_N156_wire = {M0[117], M0[137], M0[351], M0[373], M0[399], M0[547], M0[551], M0[697]};
ens0_layer0_N156 ens0_layer0_N156_inst (.M0(ens0_layer0_N156_wire), .M1(M1[156:156]));

wire [7:0] ens0_layer0_N157_wire = {M0[130], M0[191], M0[379], M0[416], M0[437], M0[712], M0[768], M0[774]};
ens0_layer0_N157 ens0_layer0_N157_inst (.M0(ens0_layer0_N157_wire), .M1(M1[157:157]));

wire [7:0] ens0_layer0_N158_wire = {M0[60], M0[79], M0[342], M0[444], M0[587], M0[639], M0[715], M0[753]};
ens0_layer0_N158 ens0_layer0_N158_inst (.M0(ens0_layer0_N158_wire), .M1(M1[158:158]));

wire [7:0] ens0_layer0_N159_wire = {M0[62], M0[339], M0[354], M0[618], M0[646], M0[652], M0[705], M0[775]};
ens0_layer0_N159 ens0_layer0_N159_inst (.M0(ens0_layer0_N159_wire), .M1(M1[159:159]));

wire [7:0] ens0_layer0_N160_wire = {M0[97], M0[195], M0[333], M0[363], M0[423], M0[524], M0[535], M0[779]};
ens0_layer0_N160 ens0_layer0_N160_inst (.M0(ens0_layer0_N160_wire), .M1(M1[160:160]));

wire [7:0] ens0_layer0_N161_wire = {M0[21], M0[108], M0[237], M0[243], M0[402], M0[589], M0[626], M0[763]};
ens0_layer0_N161 ens0_layer0_N161_inst (.M0(ens0_layer0_N161_wire), .M1(M1[161:161]));

wire [7:0] ens0_layer0_N162_wire = {M0[13], M0[72], M0[601], M0[642], M0[644], M0[727], M0[728], M0[732]};
ens0_layer0_N162 ens0_layer0_N162_inst (.M0(ens0_layer0_N162_wire), .M1(M1[162:162]));

wire [7:0] ens0_layer0_N163_wire = {M0[197], M0[228], M0[445], M0[586], M0[631], M0[684], M0[736], M0[766]};
ens0_layer0_N163 ens0_layer0_N163_inst (.M0(ens0_layer0_N163_wire), .M1(M1[163:163]));

wire [7:0] ens0_layer0_N164_wire = {M0[122], M0[196], M0[415], M0[501], M0[552], M0[579], M0[619], M0[755]};
ens0_layer0_N164 ens0_layer0_N164_inst (.M0(ens0_layer0_N164_wire), .M1(M1[164:164]));

wire [7:0] ens0_layer0_N165_wire = {M0[22], M0[289], M0[296], M0[421], M0[487], M0[600], M0[637], M0[646]};
ens0_layer0_N165 ens0_layer0_N165_inst (.M0(ens0_layer0_N165_wire), .M1(M1[165:165]));

wire [7:0] ens0_layer0_N166_wire = {M0[145], M0[170], M0[407], M0[490], M0[536], M0[642], M0[701], M0[748]};
ens0_layer0_N166 ens0_layer0_N166_inst (.M0(ens0_layer0_N166_wire), .M1(M1[166:166]));

wire [7:0] ens0_layer0_N167_wire = {M0[61], M0[214], M0[240], M0[245], M0[283], M0[518], M0[526], M0[779]};
ens0_layer0_N167 ens0_layer0_N167_inst (.M0(ens0_layer0_N167_wire), .M1(M1[167:167]));

wire [7:0] ens0_layer0_N168_wire = {M0[3], M0[10], M0[258], M0[369], M0[380], M0[570], M0[599], M0[696]};
ens0_layer0_N168 ens0_layer0_N168_inst (.M0(ens0_layer0_N168_wire), .M1(M1[168:168]));

wire [7:0] ens0_layer0_N169_wire = {M0[64], M0[152], M0[294], M0[297], M0[366], M0[442], M0[528], M0[599]};
ens0_layer0_N169 ens0_layer0_N169_inst (.M0(ens0_layer0_N169_wire), .M1(M1[169:169]));

wire [7:0] ens0_layer0_N170_wire = {M0[9], M0[58], M0[201], M0[221], M0[291], M0[423], M0[495], M0[509]};
ens0_layer0_N170 ens0_layer0_N170_inst (.M0(ens0_layer0_N170_wire), .M1(M1[170:170]));

wire [7:0] ens0_layer0_N171_wire = {M0[7], M0[93], M0[229], M0[545], M0[559], M0[660], M0[686], M0[705]};
ens0_layer0_N171 ens0_layer0_N171_inst (.M0(ens0_layer0_N171_wire), .M1(M1[171:171]));

wire [7:0] ens0_layer0_N172_wire = {M0[45], M0[101], M0[114], M0[277], M0[701], M0[740], M0[755], M0[762]};
ens0_layer0_N172 ens0_layer0_N172_inst (.M0(ens0_layer0_N172_wire), .M1(M1[172:172]));

wire [7:0] ens0_layer0_N173_wire = {M0[91], M0[110], M0[181], M0[340], M0[437], M0[502], M0[518], M0[692]};
ens0_layer0_N173 ens0_layer0_N173_inst (.M0(ens0_layer0_N173_wire), .M1(M1[173:173]));

wire [7:0] ens0_layer0_N174_wire = {M0[62], M0[180], M0[230], M0[285], M0[554], M0[597], M0[697], M0[731]};
ens0_layer0_N174 ens0_layer0_N174_inst (.M0(ens0_layer0_N174_wire), .M1(M1[174:174]));

wire [7:0] ens0_layer0_N175_wire = {M0[30], M0[41], M0[313], M0[413], M0[470], M0[503], M0[709], M0[735]};
ens0_layer0_N175 ens0_layer0_N175_inst (.M0(ens0_layer0_N175_wire), .M1(M1[175:175]));

wire [7:0] ens0_layer0_N176_wire = {M0[86], M0[95], M0[97], M0[389], M0[402], M0[403], M0[767], M0[775]};
ens0_layer0_N176 ens0_layer0_N176_inst (.M0(ens0_layer0_N176_wire), .M1(M1[176:176]));

wire [7:0] ens0_layer0_N177_wire = {M0[58], M0[99], M0[152], M0[205], M0[318], M0[373], M0[414], M0[608]};
ens0_layer0_N177 ens0_layer0_N177_inst (.M0(ens0_layer0_N177_wire), .M1(M1[177:177]));

wire [7:0] ens0_layer0_N178_wire = {M0[24], M0[44], M0[118], M0[185], M0[211], M0[447], M0[462], M0[748]};
ens0_layer0_N178 ens0_layer0_N178_inst (.M0(ens0_layer0_N178_wire), .M1(M1[178:178]));

wire [7:0] ens0_layer0_N179_wire = {M0[16], M0[40], M0[254], M0[291], M0[397], M0[527], M0[541], M0[675]};
ens0_layer0_N179 ens0_layer0_N179_inst (.M0(ens0_layer0_N179_wire), .M1(M1[179:179]));

wire [7:0] ens0_layer0_N180_wire = {M0[57], M0[415], M0[545], M0[572], M0[608], M0[660], M0[748], M0[755]};
ens0_layer0_N180 ens0_layer0_N180_inst (.M0(ens0_layer0_N180_wire), .M1(M1[180:180]));

wire [7:0] ens0_layer0_N181_wire = {M0[401], M0[421], M0[498], M0[499], M0[544], M0[587], M0[619], M0[666]};
ens0_layer0_N181 ens0_layer0_N181_inst (.M0(ens0_layer0_N181_wire), .M1(M1[181:181]));

wire [7:0] ens0_layer0_N182_wire = {M0[39], M0[239], M0[324], M0[344], M0[413], M0[444], M0[472], M0[566]};
ens0_layer0_N182 ens0_layer0_N182_inst (.M0(ens0_layer0_N182_wire), .M1(M1[182:182]));

wire [7:0] ens0_layer0_N183_wire = {M0[280], M0[308], M0[444], M0[480], M0[530], M0[649], M0[661], M0[781]};
ens0_layer0_N183 ens0_layer0_N183_inst (.M0(ens0_layer0_N183_wire), .M1(M1[183:183]));

wire [7:0] ens0_layer0_N184_wire = {M0[18], M0[187], M0[251], M0[268], M0[283], M0[493], M0[600], M0[640]};
ens0_layer0_N184 ens0_layer0_N184_inst (.M0(ens0_layer0_N184_wire), .M1(M1[184:184]));

wire [7:0] ens0_layer0_N185_wire = {M0[49], M0[58], M0[76], M0[121], M0[180], M0[493], M0[510], M0[634]};
ens0_layer0_N185 ens0_layer0_N185_inst (.M0(ens0_layer0_N185_wire), .M1(M1[185:185]));

wire [7:0] ens0_layer0_N186_wire = {M0[116], M0[190], M0[251], M0[669], M0[734], M0[744], M0[750], M0[776]};
ens0_layer0_N186 ens0_layer0_N186_inst (.M0(ens0_layer0_N186_wire), .M1(M1[186:186]));

wire [7:0] ens0_layer0_N187_wire = {M0[41], M0[197], M0[353], M0[505], M0[536], M0[595], M0[719], M0[729]};
ens0_layer0_N187 ens0_layer0_N187_inst (.M0(ens0_layer0_N187_wire), .M1(M1[187:187]));

wire [7:0] ens0_layer0_N188_wire = {M0[37], M0[159], M0[439], M0[474], M0[518], M0[537], M0[639], M0[775]};
ens0_layer0_N188 ens0_layer0_N188_inst (.M0(ens0_layer0_N188_wire), .M1(M1[188:188]));

wire [7:0] ens0_layer0_N189_wire = {M0[296], M0[320], M0[385], M0[458], M0[603], M0[696], M0[716], M0[748]};
ens0_layer0_N189 ens0_layer0_N189_inst (.M0(ens0_layer0_N189_wire), .M1(M1[189:189]));

wire [7:0] ens0_layer0_N190_wire = {M0[126], M0[220], M0[340], M0[345], M0[348], M0[626], M0[655], M0[767]};
ens0_layer0_N190 ens0_layer0_N190_inst (.M0(ens0_layer0_N190_wire), .M1(M1[190:190]));

wire [7:0] ens0_layer0_N191_wire = {M0[18], M0[85], M0[94], M0[99], M0[166], M0[264], M0[592], M0[703]};
ens0_layer0_N191 ens0_layer0_N191_inst (.M0(ens0_layer0_N191_wire), .M1(M1[191:191]));

wire [7:0] ens0_layer0_N192_wire = {M0[55], M0[98], M0[206], M0[235], M0[331], M0[460], M0[586], M0[687]};
ens0_layer0_N192 ens0_layer0_N192_inst (.M0(ens0_layer0_N192_wire), .M1(M1[192:192]));

wire [7:0] ens0_layer0_N193_wire = {M0[156], M0[383], M0[438], M0[451], M0[466], M0[490], M0[555], M0[581]};
ens0_layer0_N193 ens0_layer0_N193_inst (.M0(ens0_layer0_N193_wire), .M1(M1[193:193]));

wire [7:0] ens0_layer0_N194_wire = {M0[41], M0[126], M0[569], M0[601], M0[623], M0[625], M0[708], M0[751]};
ens0_layer0_N194 ens0_layer0_N194_inst (.M0(ens0_layer0_N194_wire), .M1(M1[194:194]));

wire [7:0] ens0_layer0_N195_wire = {M0[14], M0[170], M0[226], M0[243], M0[310], M0[312], M0[485], M0[758]};
ens0_layer0_N195 ens0_layer0_N195_inst (.M0(ens0_layer0_N195_wire), .M1(M1[195:195]));

wire [7:0] ens0_layer0_N196_wire = {M0[125], M0[143], M0[196], M0[273], M0[505], M0[522], M0[669], M0[709]};
ens0_layer0_N196 ens0_layer0_N196_inst (.M0(ens0_layer0_N196_wire), .M1(M1[196:196]));

wire [7:0] ens0_layer0_N197_wire = {M0[104], M0[258], M0[331], M0[441], M0[490], M0[578], M0[704], M0[770]};
ens0_layer0_N197 ens0_layer0_N197_inst (.M0(ens0_layer0_N197_wire), .M1(M1[197:197]));

wire [7:0] ens0_layer0_N198_wire = {M0[159], M0[236], M0[393], M0[396], M0[518], M0[634], M0[694], M0[702]};
ens0_layer0_N198 ens0_layer0_N198_inst (.M0(ens0_layer0_N198_wire), .M1(M1[198:198]));

wire [7:0] ens0_layer0_N199_wire = {M0[88], M0[260], M0[282], M0[394], M0[462], M0[533], M0[638], M0[639]};
ens0_layer0_N199 ens0_layer0_N199_inst (.M0(ens0_layer0_N199_wire), .M1(M1[199:199]));

wire [7:0] ens0_layer0_N200_wire = {M0[26], M0[124], M0[225], M0[275], M0[376], M0[597], M0[650], M0[752]};
ens0_layer0_N200 ens0_layer0_N200_inst (.M0(ens0_layer0_N200_wire), .M1(M1[200:200]));

wire [7:0] ens0_layer0_N201_wire = {M0[14], M0[175], M0[251], M0[308], M0[326], M0[377], M0[578], M0[775]};
ens0_layer0_N201 ens0_layer0_N201_inst (.M0(ens0_layer0_N201_wire), .M1(M1[201:201]));

wire [7:0] ens0_layer0_N202_wire = {M0[26], M0[116], M0[156], M0[161], M0[218], M0[449], M0[709], M0[714]};
ens0_layer0_N202 ens0_layer0_N202_inst (.M0(ens0_layer0_N202_wire), .M1(M1[202:202]));

wire [7:0] ens0_layer0_N203_wire = {M0[19], M0[53], M0[278], M0[342], M0[611], M0[655], M0[680], M0[771]};
ens0_layer0_N203 ens0_layer0_N203_inst (.M0(ens0_layer0_N203_wire), .M1(M1[203:203]));

wire [7:0] ens0_layer0_N204_wire = {M0[77], M0[295], M0[388], M0[417], M0[513], M0[523], M0[678], M0[719]};
ens0_layer0_N204 ens0_layer0_N204_inst (.M0(ens0_layer0_N204_wire), .M1(M1[204:204]));

wire [7:0] ens0_layer0_N205_wire = {M0[7], M0[203], M0[206], M0[438], M0[454], M0[568], M0[584], M0[672]};
ens0_layer0_N205 ens0_layer0_N205_inst (.M0(ens0_layer0_N205_wire), .M1(M1[205:205]));

wire [7:0] ens0_layer0_N206_wire = {M0[48], M0[105], M0[117], M0[213], M0[324], M0[452], M0[686], M0[708]};
ens0_layer0_N206 ens0_layer0_N206_inst (.M0(ens0_layer0_N206_wire), .M1(M1[206:206]));

wire [7:0] ens0_layer0_N207_wire = {M0[150], M0[216], M0[531], M0[660], M0[692], M0[708], M0[759], M0[781]};
ens0_layer0_N207 ens0_layer0_N207_inst (.M0(ens0_layer0_N207_wire), .M1(M1[207:207]));

wire [7:0] ens0_layer0_N208_wire = {M0[113], M0[196], M0[407], M0[486], M0[533], M0[609], M0[732], M0[770]};
ens0_layer0_N208 ens0_layer0_N208_inst (.M0(ens0_layer0_N208_wire), .M1(M1[208:208]));

wire [7:0] ens0_layer0_N209_wire = {M0[26], M0[70], M0[168], M0[173], M0[440], M0[521], M0[572], M0[593]};
ens0_layer0_N209 ens0_layer0_N209_inst (.M0(ens0_layer0_N209_wire), .M1(M1[209:209]));

wire [7:0] ens0_layer0_N210_wire = {M0[73], M0[139], M0[201], M0[223], M0[243], M0[329], M0[349], M0[764]};
ens0_layer0_N210 ens0_layer0_N210_inst (.M0(ens0_layer0_N210_wire), .M1(M1[210:210]));

wire [7:0] ens0_layer0_N211_wire = {M0[84], M0[146], M0[171], M0[205], M0[262], M0[479], M0[611], M0[751]};
ens0_layer0_N211 ens0_layer0_N211_inst (.M0(ens0_layer0_N211_wire), .M1(M1[211:211]));

wire [7:0] ens0_layer0_N212_wire = {M0[58], M0[200], M0[341], M0[520], M0[594], M0[670], M0[703], M0[729]};
ens0_layer0_N212 ens0_layer0_N212_inst (.M0(ens0_layer0_N212_wire), .M1(M1[212:212]));

wire [7:0] ens0_layer0_N213_wire = {M0[56], M0[77], M0[137], M0[273], M0[322], M0[339], M0[734], M0[764]};
ens0_layer0_N213 ens0_layer0_N213_inst (.M0(ens0_layer0_N213_wire), .M1(M1[213:213]));

wire [7:0] ens0_layer0_N214_wire = {M0[129], M0[236], M0[255], M0[283], M0[406], M0[432], M0[515], M0[622]};
ens0_layer0_N214 ens0_layer0_N214_inst (.M0(ens0_layer0_N214_wire), .M1(M1[214:214]));

wire [7:0] ens0_layer0_N215_wire = {M0[11], M0[100], M0[109], M0[198], M0[239], M0[349], M0[571], M0[732]};
ens0_layer0_N215 ens0_layer0_N215_inst (.M0(ens0_layer0_N215_wire), .M1(M1[215:215]));

wire [7:0] ens0_layer0_N216_wire = {M0[106], M0[125], M0[126], M0[388], M0[552], M0[563], M0[743], M0[756]};
ens0_layer0_N216 ens0_layer0_N216_inst (.M0(ens0_layer0_N216_wire), .M1(M1[216:216]));

wire [7:0] ens0_layer0_N217_wire = {M0[123], M0[144], M0[355], M0[363], M0[553], M0[618], M0[696], M0[716]};
ens0_layer0_N217 ens0_layer0_N217_inst (.M0(ens0_layer0_N217_wire), .M1(M1[217:217]));

wire [7:0] ens0_layer0_N218_wire = {M0[2], M0[43], M0[101], M0[189], M0[211], M0[522], M0[555], M0[775]};
ens0_layer0_N218 ens0_layer0_N218_inst (.M0(ens0_layer0_N218_wire), .M1(M1[218:218]));

wire [7:0] ens0_layer0_N219_wire = {M0[72], M0[355], M0[476], M0[542], M0[549], M0[680], M0[694], M0[775]};
ens0_layer0_N219 ens0_layer0_N219_inst (.M0(ens0_layer0_N219_wire), .M1(M1[219:219]));

wire [7:0] ens0_layer0_N220_wire = {M0[74], M0[160], M0[209], M0[263], M0[315], M0[522], M0[544], M0[718]};
ens0_layer0_N220 ens0_layer0_N220_inst (.M0(ens0_layer0_N220_wire), .M1(M1[220:220]));

wire [7:0] ens0_layer0_N221_wire = {M0[314], M0[379], M0[539], M0[580], M0[609], M0[648], M0[722], M0[740]};
ens0_layer0_N221 ens0_layer0_N221_inst (.M0(ens0_layer0_N221_wire), .M1(M1[221:221]));

wire [7:0] ens0_layer0_N222_wire = {M0[32], M0[70], M0[158], M0[358], M0[406], M0[518], M0[549], M0[594]};
ens0_layer0_N222 ens0_layer0_N222_inst (.M0(ens0_layer0_N222_wire), .M1(M1[222:222]));

wire [7:0] ens0_layer0_N223_wire = {M0[1], M0[261], M0[458], M0[490], M0[555], M0[583], M0[683], M0[759]};
ens0_layer0_N223 ens0_layer0_N223_inst (.M0(ens0_layer0_N223_wire), .M1(M1[223:223]));

wire [7:0] ens0_layer0_N224_wire = {M0[20], M0[169], M0[183], M0[277], M0[289], M0[524], M0[547], M0[769]};
ens0_layer0_N224 ens0_layer0_N224_inst (.M0(ens0_layer0_N224_wire), .M1(M1[224:224]));

wire [7:0] ens0_layer0_N225_wire = {M0[42], M0[276], M0[313], M0[346], M0[543], M0[735], M0[751], M0[768]};
ens0_layer0_N225 ens0_layer0_N225_inst (.M0(ens0_layer0_N225_wire), .M1(M1[225:225]));

wire [7:0] ens0_layer0_N226_wire = {M0[61], M0[67], M0[169], M0[199], M0[298], M0[359], M0[686], M0[698]};
ens0_layer0_N226 ens0_layer0_N226_inst (.M0(ens0_layer0_N226_wire), .M1(M1[226:226]));

wire [7:0] ens0_layer0_N227_wire = {M0[17], M0[127], M0[207], M0[401], M0[522], M0[546], M0[659], M0[753]};
ens0_layer0_N227 ens0_layer0_N227_inst (.M0(ens0_layer0_N227_wire), .M1(M1[227:227]));

wire [7:0] ens0_layer0_N228_wire = {M0[75], M0[80], M0[212], M0[255], M0[365], M0[499], M0[516], M0[635]};
ens0_layer0_N228 ens0_layer0_N228_inst (.M0(ens0_layer0_N228_wire), .M1(M1[228:228]));

wire [7:0] ens0_layer0_N229_wire = {M0[121], M0[217], M0[271], M0[359], M0[543], M0[670], M0[717], M0[744]};
ens0_layer0_N229 ens0_layer0_N229_inst (.M0(ens0_layer0_N229_wire), .M1(M1[229:229]));

wire [7:0] ens0_layer0_N230_wire = {M0[26], M0[30], M0[54], M0[514], M0[574], M0[589], M0[735], M0[762]};
ens0_layer0_N230 ens0_layer0_N230_inst (.M0(ens0_layer0_N230_wire), .M1(M1[230:230]));

wire [7:0] ens0_layer0_N231_wire = {M0[9], M0[50], M0[246], M0[264], M0[402], M0[677], M0[771], M0[776]};
ens0_layer0_N231 ens0_layer0_N231_inst (.M0(ens0_layer0_N231_wire), .M1(M1[231:231]));

wire [7:0] ens0_layer0_N232_wire = {M0[63], M0[99], M0[297], M0[462], M0[482], M0[508], M0[626], M0[724]};
ens0_layer0_N232 ens0_layer0_N232_inst (.M0(ens0_layer0_N232_wire), .M1(M1[232:232]));

wire [7:0] ens0_layer0_N233_wire = {M0[153], M0[216], M0[259], M0[392], M0[397], M0[579], M0[652], M0[765]};
ens0_layer0_N233 ens0_layer0_N233_inst (.M0(ens0_layer0_N233_wire), .M1(M1[233:233]));

wire [7:0] ens0_layer0_N234_wire = {M0[28], M0[34], M0[223], M0[330], M0[381], M0[480], M0[492], M0[732]};
ens0_layer0_N234 ens0_layer0_N234_inst (.M0(ens0_layer0_N234_wire), .M1(M1[234:234]));

wire [7:0] ens0_layer0_N235_wire = {M0[286], M0[318], M0[320], M0[366], M0[456], M0[533], M0[654], M0[783]};
ens0_layer0_N235 ens0_layer0_N235_inst (.M0(ens0_layer0_N235_wire), .M1(M1[235:235]));

wire [7:0] ens0_layer0_N236_wire = {M0[97], M0[121], M0[423], M0[491], M0[564], M0[683], M0[737], M0[753]};
ens0_layer0_N236 ens0_layer0_N236_inst (.M0(ens0_layer0_N236_wire), .M1(M1[236:236]));

wire [7:0] ens0_layer0_N237_wire = {M0[37], M0[139], M0[368], M0[474], M0[477], M0[480], M0[620], M0[756]};
ens0_layer0_N237 ens0_layer0_N237_inst (.M0(ens0_layer0_N237_wire), .M1(M1[237:237]));

wire [7:0] ens0_layer0_N238_wire = {M0[38], M0[52], M0[211], M0[228], M0[346], M0[493], M0[558], M0[715]};
ens0_layer0_N238 ens0_layer0_N238_inst (.M0(ens0_layer0_N238_wire), .M1(M1[238:238]));

wire [7:0] ens0_layer0_N239_wire = {M0[16], M0[31], M0[152], M0[160], M0[188], M0[327], M0[480], M0[733]};
ens0_layer0_N239 ens0_layer0_N239_inst (.M0(ens0_layer0_N239_wire), .M1(M1[239:239]));

wire [7:0] ens0_layer0_N240_wire = {M0[67], M0[128], M0[143], M0[529], M0[562], M0[564], M0[661], M0[755]};
ens0_layer0_N240 ens0_layer0_N240_inst (.M0(ens0_layer0_N240_wire), .M1(M1[240:240]));

wire [7:0] ens0_layer0_N241_wire = {M0[4], M0[213], M0[305], M0[332], M0[398], M0[638], M0[721], M0[728]};
ens0_layer0_N241 ens0_layer0_N241_inst (.M0(ens0_layer0_N241_wire), .M1(M1[241:241]));

wire [7:0] ens0_layer0_N242_wire = {M0[21], M0[34], M0[280], M0[347], M0[351], M0[510], M0[572], M0[596]};
ens0_layer0_N242 ens0_layer0_N242_inst (.M0(ens0_layer0_N242_wire), .M1(M1[242:242]));

wire [7:0] ens0_layer0_N243_wire = {M0[27], M0[230], M0[262], M0[380], M0[406], M0[425], M0[729], M0[782]};
ens0_layer0_N243 ens0_layer0_N243_inst (.M0(ens0_layer0_N243_wire), .M1(M1[243:243]));

wire [7:0] ens0_layer0_N244_wire = {M0[60], M0[209], M0[213], M0[346], M0[397], M0[559], M0[592], M0[639]};
ens0_layer0_N244 ens0_layer0_N244_inst (.M0(ens0_layer0_N244_wire), .M1(M1[244:244]));

wire [7:0] ens0_layer0_N245_wire = {M0[16], M0[327], M0[399], M0[424], M0[448], M0[497], M0[593], M0[731]};
ens0_layer0_N245 ens0_layer0_N245_inst (.M0(ens0_layer0_N245_wire), .M1(M1[245:245]));

wire [7:0] ens0_layer0_N246_wire = {M0[92], M0[162], M0[366], M0[427], M0[495], M0[640], M0[645], M0[744]};
ens0_layer0_N246 ens0_layer0_N246_inst (.M0(ens0_layer0_N246_wire), .M1(M1[246:246]));

wire [7:0] ens0_layer0_N247_wire = {M0[424], M0[466], M0[505], M0[587], M0[588], M0[613], M0[624], M0[748]};
ens0_layer0_N247 ens0_layer0_N247_inst (.M0(ens0_layer0_N247_wire), .M1(M1[247:247]));

wire [7:0] ens0_layer0_N248_wire = {M0[66], M0[203], M0[217], M0[253], M0[352], M0[641], M0[651], M0[712]};
ens0_layer0_N248 ens0_layer0_N248_inst (.M0(ens0_layer0_N248_wire), .M1(M1[248:248]));

wire [7:0] ens0_layer0_N249_wire = {M0[109], M0[125], M0[165], M0[187], M0[315], M0[336], M0[388], M0[712]};
ens0_layer0_N249 ens0_layer0_N249_inst (.M0(ens0_layer0_N249_wire), .M1(M1[249:249]));

wire [7:0] ens0_layer0_N250_wire = {M0[391], M0[411], M0[464], M0[469], M0[616], M0[620], M0[653], M0[735]};
ens0_layer0_N250 ens0_layer0_N250_inst (.M0(ens0_layer0_N250_wire), .M1(M1[250:250]));

wire [7:0] ens0_layer0_N251_wire = {M0[37], M0[167], M0[298], M0[304], M0[342], M0[377], M0[690], M0[744]};
ens0_layer0_N251 ens0_layer0_N251_inst (.M0(ens0_layer0_N251_wire), .M1(M1[251:251]));

wire [7:0] ens0_layer0_N252_wire = {M0[67], M0[104], M0[125], M0[340], M0[476], M0[519], M0[655], M0[703]};
ens0_layer0_N252 ens0_layer0_N252_inst (.M0(ens0_layer0_N252_wire), .M1(M1[252:252]));

wire [7:0] ens0_layer0_N253_wire = {M0[90], M0[153], M0[423], M0[442], M0[444], M0[563], M0[693], M0[769]};
ens0_layer0_N253 ens0_layer0_N253_inst (.M0(ens0_layer0_N253_wire), .M1(M1[253:253]));

wire [7:0] ens0_layer0_N254_wire = {M0[145], M0[166], M0[238], M0[271], M0[411], M0[482], M0[588], M0[782]};
ens0_layer0_N254 ens0_layer0_N254_inst (.M0(ens0_layer0_N254_wire), .M1(M1[254:254]));

wire [7:0] ens0_layer0_N255_wire = {M0[193], M0[208], M0[233], M0[293], M0[414], M0[458], M0[594], M0[759]};
ens0_layer0_N255 ens0_layer0_N255_inst (.M0(ens0_layer0_N255_wire), .M1(M1[255:255]));

wire [7:0] ens0_layer0_N256_wire = {M0[66], M0[305], M0[345], M0[365], M0[366], M0[432], M0[496], M0[554]};
ens0_layer0_N256 ens0_layer0_N256_inst (.M0(ens0_layer0_N256_wire), .M1(M1[256:256]));

wire [7:0] ens0_layer0_N257_wire = {M0[23], M0[115], M0[143], M0[152], M0[177], M0[178], M0[314], M0[343]};
ens0_layer0_N257 ens0_layer0_N257_inst (.M0(ens0_layer0_N257_wire), .M1(M1[257:257]));

wire [7:0] ens0_layer0_N258_wire = {M0[45], M0[89], M0[140], M0[258], M0[331], M0[356], M0[599], M0[613]};
ens0_layer0_N258 ens0_layer0_N258_inst (.M0(ens0_layer0_N258_wire), .M1(M1[258:258]));

wire [7:0] ens0_layer0_N259_wire = {M0[100], M0[132], M0[180], M0[202], M0[266], M0[320], M0[545], M0[602]};
ens0_layer0_N259 ens0_layer0_N259_inst (.M0(ens0_layer0_N259_wire), .M1(M1[259:259]));

wire [7:0] ens0_layer0_N260_wire = {M0[135], M0[237], M0[339], M0[347], M0[398], M0[498], M0[655], M0[701]};
ens0_layer0_N260 ens0_layer0_N260_inst (.M0(ens0_layer0_N260_wire), .M1(M1[260:260]));

wire [7:0] ens0_layer0_N261_wire = {M0[189], M0[240], M0[301], M0[373], M0[428], M0[490], M0[582], M0[702]};
ens0_layer0_N261 ens0_layer0_N261_inst (.M0(ens0_layer0_N261_wire), .M1(M1[261:261]));

wire [7:0] ens0_layer0_N262_wire = {M0[40], M0[70], M0[118], M0[130], M0[265], M0[306], M0[426], M0[494]};
ens0_layer0_N262 ens0_layer0_N262_inst (.M0(ens0_layer0_N262_wire), .M1(M1[262:262]));

wire [7:0] ens0_layer0_N263_wire = {M0[137], M0[222], M0[289], M0[304], M0[319], M0[352], M0[425], M0[474]};
ens0_layer0_N263 ens0_layer0_N263_inst (.M0(ens0_layer0_N263_wire), .M1(M1[263:263]));

wire [7:0] ens0_layer0_N264_wire = {M0[110], M0[222], M0[252], M0[259], M0[378], M0[448], M0[600], M0[741]};
ens0_layer0_N264 ens0_layer0_N264_inst (.M0(ens0_layer0_N264_wire), .M1(M1[264:264]));

wire [7:0] ens0_layer0_N265_wire = {M0[262], M0[315], M0[331], M0[393], M0[447], M0[480], M0[521], M0[547]};
ens0_layer0_N265 ens0_layer0_N265_inst (.M0(ens0_layer0_N265_wire), .M1(M1[265:265]));

wire [7:0] ens0_layer0_N266_wire = {M0[51], M0[107], M0[233], M0[336], M0[422], M0[435], M0[547], M0[646]};
ens0_layer0_N266 ens0_layer0_N266_inst (.M0(ens0_layer0_N266_wire), .M1(M1[266:266]));

wire [7:0] ens0_layer0_N267_wire = {M0[3], M0[19], M0[60], M0[313], M0[574], M0[606], M0[614], M0[731]};
ens0_layer0_N267 ens0_layer0_N267_inst (.M0(ens0_layer0_N267_wire), .M1(M1[267:267]));

wire [7:0] ens0_layer0_N268_wire = {M0[98], M0[139], M0[164], M0[214], M0[393], M0[396], M0[503], M0[624]};
ens0_layer0_N268 ens0_layer0_N268_inst (.M0(ens0_layer0_N268_wire), .M1(M1[268:268]));

wire [7:0] ens0_layer0_N269_wire = {M0[96], M0[155], M0[426], M0[515], M0[665], M0[696], M0[765], M0[783]};
ens0_layer0_N269 ens0_layer0_N269_inst (.M0(ens0_layer0_N269_wire), .M1(M1[269:269]));

wire [7:0] ens0_layer0_N270_wire = {M0[21], M0[26], M0[61], M0[77], M0[304], M0[514], M0[662], M0[673]};
ens0_layer0_N270 ens0_layer0_N270_inst (.M0(ens0_layer0_N270_wire), .M1(M1[270:270]));

wire [7:0] ens0_layer0_N271_wire = {M0[101], M0[222], M0[224], M0[505], M0[580], M0[651], M0[707], M0[770]};
ens0_layer0_N271 ens0_layer0_N271_inst (.M0(ens0_layer0_N271_wire), .M1(M1[271:271]));

wire [7:0] ens0_layer0_N272_wire = {M0[264], M0[326], M0[419], M0[550], M0[576], M0[618], M0[620], M0[769]};
ens0_layer0_N272 ens0_layer0_N272_inst (.M0(ens0_layer0_N272_wire), .M1(M1[272:272]));

wire [7:0] ens0_layer0_N273_wire = {M0[241], M0[370], M0[447], M0[519], M0[541], M0[592], M0[633], M0[674]};
ens0_layer0_N273 ens0_layer0_N273_inst (.M0(ens0_layer0_N273_wire), .M1(M1[273:273]));

wire [7:0] ens0_layer0_N274_wire = {M0[141], M0[213], M0[224], M0[359], M0[582], M0[613], M0[653], M0[722]};
ens0_layer0_N274 ens0_layer0_N274_inst (.M0(ens0_layer0_N274_wire), .M1(M1[274:274]));

wire [7:0] ens0_layer0_N275_wire = {M0[69], M0[179], M0[273], M0[337], M0[338], M0[450], M0[478], M0[766]};
ens0_layer0_N275 ens0_layer0_N275_inst (.M0(ens0_layer0_N275_wire), .M1(M1[275:275]));

wire [7:0] ens0_layer0_N276_wire = {M0[30], M0[59], M0[90], M0[273], M0[369], M0[421], M0[660], M0[748]};
ens0_layer0_N276 ens0_layer0_N276_inst (.M0(ens0_layer0_N276_wire), .M1(M1[276:276]));

wire [7:0] ens0_layer0_N277_wire = {M0[16], M0[127], M0[176], M0[242], M0[334], M0[397], M0[399], M0[640]};
ens0_layer0_N277 ens0_layer0_N277_inst (.M0(ens0_layer0_N277_wire), .M1(M1[277:277]));

wire [7:0] ens0_layer0_N278_wire = {M0[68], M0[119], M0[140], M0[286], M0[392], M0[395], M0[625], M0[693]};
ens0_layer0_N278 ens0_layer0_N278_inst (.M0(ens0_layer0_N278_wire), .M1(M1[278:278]));

wire [7:0] ens0_layer0_N279_wire = {M0[35], M0[68], M0[90], M0[132], M0[143], M0[254], M0[463], M0[732]};
ens0_layer0_N279 ens0_layer0_N279_inst (.M0(ens0_layer0_N279_wire), .M1(M1[279:279]));

wire [7:0] ens0_layer0_N280_wire = {M0[183], M0[261], M0[310], M0[396], M0[463], M0[499], M0[556], M0[639]};
ens0_layer0_N280 ens0_layer0_N280_inst (.M0(ens0_layer0_N280_wire), .M1(M1[280:280]));

wire [7:0] ens0_layer0_N281_wire = {M0[54], M0[173], M0[193], M0[416], M0[468], M0[641], M0[645], M0[659]};
ens0_layer0_N281 ens0_layer0_N281_inst (.M0(ens0_layer0_N281_wire), .M1(M1[281:281]));

wire [7:0] ens0_layer0_N282_wire = {M0[69], M0[143], M0[292], M0[425], M0[477], M0[496], M0[526], M0[702]};
ens0_layer0_N282 ens0_layer0_N282_inst (.M0(ens0_layer0_N282_wire), .M1(M1[282:282]));

wire [7:0] ens0_layer0_N283_wire = {M0[23], M0[94], M0[180], M0[400], M0[517], M0[624], M0[691], M0[779]};
ens0_layer0_N283 ens0_layer0_N283_inst (.M0(ens0_layer0_N283_wire), .M1(M1[283:283]));

wire [7:0] ens0_layer0_N284_wire = {M0[175], M0[233], M0[250], M0[286], M0[321], M0[388], M0[515], M0[618]};
ens0_layer0_N284 ens0_layer0_N284_inst (.M0(ens0_layer0_N284_wire), .M1(M1[284:284]));

wire [7:0] ens0_layer0_N285_wire = {M0[0], M0[38], M0[77], M0[126], M0[179], M0[498], M0[641], M0[722]};
ens0_layer0_N285 ens0_layer0_N285_inst (.M0(ens0_layer0_N285_wire), .M1(M1[285:285]));

wire [7:0] ens0_layer0_N286_wire = {M0[47], M0[197], M0[211], M0[375], M0[453], M0[550], M0[703], M0[780]};
ens0_layer0_N286 ens0_layer0_N286_inst (.M0(ens0_layer0_N286_wire), .M1(M1[286:286]));

wire [7:0] ens0_layer0_N287_wire = {M0[23], M0[58], M0[399], M0[516], M0[635], M0[665], M0[713], M0[736]};
ens0_layer0_N287 ens0_layer0_N287_inst (.M0(ens0_layer0_N287_wire), .M1(M1[287:287]));

wire [7:0] ens0_layer0_N288_wire = {M0[89], M0[288], M0[309], M0[364], M0[538], M0[604], M0[740], M0[778]};
ens0_layer0_N288 ens0_layer0_N288_inst (.M0(ens0_layer0_N288_wire), .M1(M1[288:288]));

wire [7:0] ens0_layer0_N289_wire = {M0[97], M0[187], M0[220], M0[230], M0[361], M0[387], M0[402], M0[548]};
ens0_layer0_N289 ens0_layer0_N289_inst (.M0(ens0_layer0_N289_wire), .M1(M1[289:289]));

wire [7:0] ens0_layer0_N290_wire = {M0[81], M0[160], M0[162], M0[224], M0[278], M0[345], M0[393], M0[732]};
ens0_layer0_N290 ens0_layer0_N290_inst (.M0(ens0_layer0_N290_wire), .M1(M1[290:290]));

wire [7:0] ens0_layer0_N291_wire = {M0[254], M0[345], M0[431], M0[449], M0[538], M0[575], M0[585], M0[696]};
ens0_layer0_N291 ens0_layer0_N291_inst (.M0(ens0_layer0_N291_wire), .M1(M1[291:291]));

wire [7:0] ens0_layer0_N292_wire = {M0[51], M0[101], M0[378], M0[423], M0[558], M0[576], M0[578], M0[659]};
ens0_layer0_N292 ens0_layer0_N292_inst (.M0(ens0_layer0_N292_wire), .M1(M1[292:292]));

wire [7:0] ens0_layer0_N293_wire = {M0[25], M0[80], M0[81], M0[93], M0[263], M0[527], M0[576], M0[698]};
ens0_layer0_N293 ens0_layer0_N293_inst (.M0(ens0_layer0_N293_wire), .M1(M1[293:293]));

wire [7:0] ens0_layer0_N294_wire = {M0[65], M0[294], M0[338], M0[445], M0[513], M0[601], M0[698], M0[705]};
ens0_layer0_N294 ens0_layer0_N294_inst (.M0(ens0_layer0_N294_wire), .M1(M1[294:294]));

wire [7:0] ens0_layer0_N295_wire = {M0[52], M0[388], M0[406], M0[417], M0[479], M0[497], M0[499], M0[608]};
ens0_layer0_N295 ens0_layer0_N295_inst (.M0(ens0_layer0_N295_wire), .M1(M1[295:295]));

wire [7:0] ens0_layer0_N296_wire = {M0[19], M0[56], M0[233], M0[299], M0[451], M0[465], M0[537], M0[715]};
ens0_layer0_N296 ens0_layer0_N296_inst (.M0(ens0_layer0_N296_wire), .M1(M1[296:296]));

wire [7:0] ens0_layer0_N297_wire = {M0[36], M0[144], M0[206], M0[333], M0[393], M0[562], M0[747], M0[780]};
ens0_layer0_N297 ens0_layer0_N297_inst (.M0(ens0_layer0_N297_wire), .M1(M1[297:297]));

wire [7:0] ens0_layer0_N298_wire = {M0[230], M0[324], M0[325], M0[577], M0[655], M0[660], M0[742], M0[743]};
ens0_layer0_N298 ens0_layer0_N298_inst (.M0(ens0_layer0_N298_wire), .M1(M1[298:298]));

wire [7:0] ens0_layer0_N299_wire = {M0[41], M0[213], M0[301], M0[466], M0[500], M0[546], M0[746], M0[781]};
ens0_layer0_N299 ens0_layer0_N299_inst (.M0(ens0_layer0_N299_wire), .M1(M1[299:299]));

wire [7:0] ens0_layer0_N300_wire = {M0[18], M0[58], M0[118], M0[154], M0[165], M0[417], M0[519], M0[536]};
ens0_layer0_N300 ens0_layer0_N300_inst (.M0(ens0_layer0_N300_wire), .M1(M1[300:300]));

wire [7:0] ens0_layer0_N301_wire = {M0[126], M0[141], M0[156], M0[220], M0[309], M0[477], M0[689], M0[737]};
ens0_layer0_N301 ens0_layer0_N301_inst (.M0(ens0_layer0_N301_wire), .M1(M1[301:301]));

wire [7:0] ens0_layer0_N302_wire = {M0[174], M0[187], M0[234], M0[313], M0[374], M0[479], M0[584], M0[617]};
ens0_layer0_N302 ens0_layer0_N302_inst (.M0(ens0_layer0_N302_wire), .M1(M1[302:302]));

wire [7:0] ens0_layer0_N303_wire = {M0[4], M0[84], M0[99], M0[202], M0[352], M0[368], M0[472], M0[671]};
ens0_layer0_N303 ens0_layer0_N303_inst (.M0(ens0_layer0_N303_wire), .M1(M1[303:303]));

wire [7:0] ens0_layer0_N304_wire = {M0[33], M0[241], M0[293], M0[345], M0[519], M0[633], M0[732], M0[738]};
ens0_layer0_N304 ens0_layer0_N304_inst (.M0(ens0_layer0_N304_wire), .M1(M1[304:304]));

wire [7:0] ens0_layer0_N305_wire = {M0[14], M0[40], M0[56], M0[105], M0[201], M0[345], M0[497], M0[549]};
ens0_layer0_N305 ens0_layer0_N305_inst (.M0(ens0_layer0_N305_wire), .M1(M1[305:305]));

wire [7:0] ens0_layer0_N306_wire = {M0[70], M0[199], M0[233], M0[411], M0[515], M0[638], M0[673], M0[772]};
ens0_layer0_N306 ens0_layer0_N306_inst (.M0(ens0_layer0_N306_wire), .M1(M1[306:306]));

wire [7:0] ens0_layer0_N307_wire = {M0[138], M0[496], M0[528], M0[529], M0[697], M0[714], M0[725], M0[774]};
ens0_layer0_N307 ens0_layer0_N307_inst (.M0(ens0_layer0_N307_wire), .M1(M1[307:307]));

wire [7:0] ens0_layer0_N308_wire = {M0[70], M0[100], M0[159], M0[349], M0[354], M0[455], M0[603], M0[642]};
ens0_layer0_N308 ens0_layer0_N308_inst (.M0(ens0_layer0_N308_wire), .M1(M1[308:308]));

wire [7:0] ens0_layer0_N309_wire = {M0[17], M0[42], M0[64], M0[70], M0[82], M0[357], M0[369], M0[637]};
ens0_layer0_N309 ens0_layer0_N309_inst (.M0(ens0_layer0_N309_wire), .M1(M1[309:309]));

wire [7:0] ens0_layer0_N310_wire = {M0[16], M0[130], M0[415], M0[429], M0[454], M0[601], M0[632], M0[730]};
ens0_layer0_N310 ens0_layer0_N310_inst (.M0(ens0_layer0_N310_wire), .M1(M1[310:310]));

wire [7:0] ens0_layer0_N311_wire = {M0[6], M0[34], M0[432], M0[441], M0[643], M0[700], M0[705], M0[770]};
ens0_layer0_N311 ens0_layer0_N311_inst (.M0(ens0_layer0_N311_wire), .M1(M1[311:311]));

wire [7:0] ens0_layer0_N312_wire = {M0[60], M0[224], M0[227], M0[289], M0[327], M0[359], M0[558], M0[604]};
ens0_layer0_N312 ens0_layer0_N312_inst (.M0(ens0_layer0_N312_wire), .M1(M1[312:312]));

wire [7:0] ens0_layer0_N313_wire = {M0[352], M0[365], M0[402], M0[550], M0[631], M0[660], M0[768], M0[770]};
ens0_layer0_N313 ens0_layer0_N313_inst (.M0(ens0_layer0_N313_wire), .M1(M1[313:313]));

wire [7:0] ens0_layer0_N314_wire = {M0[218], M0[347], M0[401], M0[421], M0[447], M0[489], M0[507], M0[740]};
ens0_layer0_N314 ens0_layer0_N314_inst (.M0(ens0_layer0_N314_wire), .M1(M1[314:314]));

wire [7:0] ens0_layer0_N315_wire = {M0[0], M0[82], M0[386], M0[497], M0[503], M0[578], M0[597], M0[653]};
ens0_layer0_N315 ens0_layer0_N315_inst (.M0(ens0_layer0_N315_wire), .M1(M1[315:315]));

wire [7:0] ens0_layer0_N316_wire = {M0[138], M0[336], M0[390], M0[406], M0[472], M0[506], M0[555], M0[586]};
ens0_layer0_N316 ens0_layer0_N316_inst (.M0(ens0_layer0_N316_wire), .M1(M1[316:316]));

wire [7:0] ens0_layer0_N317_wire = {M0[142], M0[179], M0[313], M0[341], M0[509], M0[627], M0[696], M0[758]};
ens0_layer0_N317 ens0_layer0_N317_inst (.M0(ens0_layer0_N317_wire), .M1(M1[317:317]));

wire [7:0] ens0_layer0_N318_wire = {M0[135], M0[159], M0[177], M0[510], M0[532], M0[575], M0[640], M0[654]};
ens0_layer0_N318 ens0_layer0_N318_inst (.M0(ens0_layer0_N318_wire), .M1(M1[318:318]));

wire [7:0] ens0_layer0_N319_wire = {M0[36], M0[210], M0[256], M0[321], M0[403], M0[680], M0[692], M0[742]};
ens0_layer0_N319 ens0_layer0_N319_inst (.M0(ens0_layer0_N319_wire), .M1(M1[319:319]));

wire [7:0] ens0_layer0_N320_wire = {M0[6], M0[200], M0[416], M0[449], M0[578], M0[605], M0[702], M0[775]};
ens0_layer0_N320 ens0_layer0_N320_inst (.M0(ens0_layer0_N320_wire), .M1(M1[320:320]));

wire [7:0] ens0_layer0_N321_wire = {M0[130], M0[313], M0[337], M0[344], M0[363], M0[456], M0[484], M0[676]};
ens0_layer0_N321 ens0_layer0_N321_inst (.M0(ens0_layer0_N321_wire), .M1(M1[321:321]));

wire [7:0] ens0_layer0_N322_wire = {M0[68], M0[372], M0[459], M0[620], M0[634], M0[651], M0[687], M0[733]};
ens0_layer0_N322 ens0_layer0_N322_inst (.M0(ens0_layer0_N322_wire), .M1(M1[322:322]));

wire [7:0] ens0_layer0_N323_wire = {M0[249], M0[379], M0[442], M0[471], M0[561], M0[576], M0[713], M0[744]};
ens0_layer0_N323 ens0_layer0_N323_inst (.M0(ens0_layer0_N323_wire), .M1(M1[323:323]));

wire [7:0] ens0_layer0_N324_wire = {M0[212], M0[326], M0[352], M0[464], M0[545], M0[589], M0[639], M0[774]};
ens0_layer0_N324 ens0_layer0_N324_inst (.M0(ens0_layer0_N324_wire), .M1(M1[324:324]));

wire [7:0] ens0_layer0_N325_wire = {M0[244], M0[266], M0[292], M0[299], M0[371], M0[498], M0[614], M0[751]};
ens0_layer0_N325 ens0_layer0_N325_inst (.M0(ens0_layer0_N325_wire), .M1(M1[325:325]));

wire [7:0] ens0_layer0_N326_wire = {M0[103], M0[140], M0[311], M0[349], M0[506], M0[611], M0[684], M0[736]};
ens0_layer0_N326 ens0_layer0_N326_inst (.M0(ens0_layer0_N326_wire), .M1(M1[326:326]));

wire [7:0] ens0_layer0_N327_wire = {M0[162], M0[299], M0[357], M0[407], M0[553], M0[634], M0[703], M0[725]};
ens0_layer0_N327 ens0_layer0_N327_inst (.M0(ens0_layer0_N327_wire), .M1(M1[327:327]));

wire [7:0] ens0_layer0_N328_wire = {M0[97], M0[270], M0[298], M0[333], M0[354], M0[355], M0[509], M0[723]};
ens0_layer0_N328 ens0_layer0_N328_inst (.M0(ens0_layer0_N328_wire), .M1(M1[328:328]));

wire [7:0] ens0_layer0_N329_wire = {M0[14], M0[138], M0[265], M0[276], M0[448], M0[474], M0[511], M0[658]};
ens0_layer0_N329 ens0_layer0_N329_inst (.M0(ens0_layer0_N329_wire), .M1(M1[329:329]));

wire [7:0] ens0_layer0_N330_wire = {M0[12], M0[75], M0[115], M0[152], M0[175], M0[227], M0[379], M0[695]};
ens0_layer0_N330 ens0_layer0_N330_inst (.M0(ens0_layer0_N330_wire), .M1(M1[330:330]));

wire [7:0] ens0_layer0_N331_wire = {M0[138], M0[165], M0[433], M0[531], M0[672], M0[673], M0[675], M0[681]};
ens0_layer0_N331 ens0_layer0_N331_inst (.M0(ens0_layer0_N331_wire), .M1(M1[331:331]));

wire [7:0] ens0_layer0_N332_wire = {M0[151], M0[161], M0[261], M0[325], M0[428], M0[483], M0[619], M0[696]};
ens0_layer0_N332 ens0_layer0_N332_inst (.M0(ens0_layer0_N332_wire), .M1(M1[332:332]));

wire [7:0] ens0_layer0_N333_wire = {M0[13], M0[25], M0[120], M0[351], M0[501], M0[509], M0[761], M0[778]};
ens0_layer0_N333 ens0_layer0_N333_inst (.M0(ens0_layer0_N333_wire), .M1(M1[333:333]));

wire [7:0] ens0_layer0_N334_wire = {M0[210], M0[241], M0[306], M0[342], M0[558], M0[612], M0[614], M0[751]};
ens0_layer0_N334 ens0_layer0_N334_inst (.M0(ens0_layer0_N334_wire), .M1(M1[334:334]));

wire [7:0] ens0_layer0_N335_wire = {M0[49], M0[83], M0[305], M0[306], M0[333], M0[560], M0[576], M0[669]};
ens0_layer0_N335 ens0_layer0_N335_inst (.M0(ens0_layer0_N335_wire), .M1(M1[335:335]));

wire [7:0] ens0_layer0_N336_wire = {M0[351], M0[558], M0[570], M0[626], M0[670], M0[714], M0[727], M0[767]};
ens0_layer0_N336 ens0_layer0_N336_inst (.M0(ens0_layer0_N336_wire), .M1(M1[336:336]));

wire [7:0] ens0_layer0_N337_wire = {M0[99], M0[105], M0[153], M0[191], M0[409], M0[531], M0[598], M0[659]};
ens0_layer0_N337 ens0_layer0_N337_inst (.M0(ens0_layer0_N337_wire), .M1(M1[337:337]));

wire [7:0] ens0_layer0_N338_wire = {M0[36], M0[113], M0[153], M0[337], M0[382], M0[532], M0[539], M0[724]};
ens0_layer0_N338 ens0_layer0_N338_inst (.M0(ens0_layer0_N338_wire), .M1(M1[338:338]));

wire [7:0] ens0_layer0_N339_wire = {M0[22], M0[34], M0[168], M0[435], M0[472], M0[608], M0[628], M0[769]};
ens0_layer0_N339 ens0_layer0_N339_inst (.M0(ens0_layer0_N339_wire), .M1(M1[339:339]));

wire [7:0] ens0_layer0_N340_wire = {M0[39], M0[85], M0[149], M0[417], M0[428], M0[486], M0[626], M0[691]};
ens0_layer0_N340 ens0_layer0_N340_inst (.M0(ens0_layer0_N340_wire), .M1(M1[340:340]));

wire [7:0] ens0_layer0_N341_wire = {M0[27], M0[62], M0[64], M0[72], M0[202], M0[494], M0[524], M0[530]};
ens0_layer0_N341 ens0_layer0_N341_inst (.M0(ens0_layer0_N341_wire), .M1(M1[341:341]));

wire [7:0] ens0_layer0_N342_wire = {M0[270], M0[397], M0[427], M0[460], M0[493], M0[627], M0[693], M0[741]};
ens0_layer0_N342 ens0_layer0_N342_inst (.M0(ens0_layer0_N342_wire), .M1(M1[342:342]));

wire [7:0] ens0_layer0_N343_wire = {M0[9], M0[103], M0[104], M0[132], M0[199], M0[630], M0[778], M0[779]};
ens0_layer0_N343 ens0_layer0_N343_inst (.M0(ens0_layer0_N343_wire), .M1(M1[343:343]));

wire [7:0] ens0_layer0_N344_wire = {M0[195], M0[196], M0[354], M0[402], M0[518], M0[538], M0[623], M0[646]};
ens0_layer0_N344 ens0_layer0_N344_inst (.M0(ens0_layer0_N344_wire), .M1(M1[344:344]));

wire [7:0] ens0_layer0_N345_wire = {M0[40], M0[193], M0[226], M0[354], M0[621], M0[625], M0[658], M0[774]};
ens0_layer0_N345 ens0_layer0_N345_inst (.M0(ens0_layer0_N345_wire), .M1(M1[345:345]));

wire [7:0] ens0_layer0_N346_wire = {M0[5], M0[114], M0[250], M0[334], M0[394], M0[549], M0[620], M0[623]};
ens0_layer0_N346 ens0_layer0_N346_inst (.M0(ens0_layer0_N346_wire), .M1(M1[346:346]));

wire [7:0] ens0_layer0_N347_wire = {M0[30], M0[37], M0[200], M0[292], M0[302], M0[370], M0[445], M0[459]};
ens0_layer0_N347 ens0_layer0_N347_inst (.M0(ens0_layer0_N347_wire), .M1(M1[347:347]));

wire [7:0] ens0_layer0_N348_wire = {M0[20], M0[107], M0[177], M0[280], M0[307], M0[360], M0[540], M0[569]};
ens0_layer0_N348 ens0_layer0_N348_inst (.M0(ens0_layer0_N348_wire), .M1(M1[348:348]));

wire [7:0] ens0_layer0_N349_wire = {M0[27], M0[28], M0[61], M0[276], M0[421], M0[587], M0[693], M0[694]};
ens0_layer0_N349 ens0_layer0_N349_inst (.M0(ens0_layer0_N349_wire), .M1(M1[349:349]));

wire [7:0] ens0_layer0_N350_wire = {M0[101], M0[250], M0[417], M0[431], M0[540], M0[565], M0[648], M0[694]};
ens0_layer0_N350 ens0_layer0_N350_inst (.M0(ens0_layer0_N350_wire), .M1(M1[350:350]));

wire [7:0] ens0_layer0_N351_wire = {M0[183], M0[212], M0[258], M0[498], M0[586], M0[656], M0[662], M0[768]};
ens0_layer0_N351 ens0_layer0_N351_inst (.M0(ens0_layer0_N351_wire), .M1(M1[351:351]));

wire [7:0] ens0_layer0_N352_wire = {M0[13], M0[90], M0[172], M0[345], M0[355], M0[384], M0[562], M0[586]};
ens0_layer0_N352 ens0_layer0_N352_inst (.M0(ens0_layer0_N352_wire), .M1(M1[352:352]));

wire [7:0] ens0_layer0_N353_wire = {M0[14], M0[23], M0[38], M0[57], M0[103], M0[406], M0[525], M0[533]};
ens0_layer0_N353 ens0_layer0_N353_inst (.M0(ens0_layer0_N353_wire), .M1(M1[353:353]));

wire [7:0] ens0_layer0_N354_wire = {M0[347], M0[416], M0[436], M0[638], M0[679], M0[696], M0[708], M0[774]};
ens0_layer0_N354 ens0_layer0_N354_inst (.M0(ens0_layer0_N354_wire), .M1(M1[354:354]));

wire [7:0] ens0_layer0_N355_wire = {M0[177], M0[245], M0[296], M0[313], M0[585], M0[601], M0[685], M0[723]};
ens0_layer0_N355 ens0_layer0_N355_inst (.M0(ens0_layer0_N355_wire), .M1(M1[355:355]));

wire [7:0] ens0_layer0_N356_wire = {M0[183], M0[223], M0[262], M0[316], M0[372], M0[525], M0[555], M0[691]};
ens0_layer0_N356 ens0_layer0_N356_inst (.M0(ens0_layer0_N356_wire), .M1(M1[356:356]));

wire [7:0] ens0_layer0_N357_wire = {M0[17], M0[292], M0[385], M0[488], M0[514], M0[618], M0[724], M0[769]};
ens0_layer0_N357 ens0_layer0_N357_inst (.M0(ens0_layer0_N357_wire), .M1(M1[357:357]));

wire [7:0] ens0_layer0_N358_wire = {M0[24], M0[26], M0[89], M0[337], M0[517], M0[608], M0[616], M0[748]};
ens0_layer0_N358 ens0_layer0_N358_inst (.M0(ens0_layer0_N358_wire), .M1(M1[358:358]));

wire [7:0] ens0_layer0_N359_wire = {M0[131], M0[285], M0[316], M0[364], M0[538], M0[681], M0[716], M0[754]};
ens0_layer0_N359 ens0_layer0_N359_inst (.M0(ens0_layer0_N359_wire), .M1(M1[359:359]));

wire [7:0] ens0_layer0_N360_wire = {M0[50], M0[236], M0[241], M0[367], M0[463], M0[547], M0[689], M0[757]};
ens0_layer0_N360 ens0_layer0_N360_inst (.M0(ens0_layer0_N360_wire), .M1(M1[360:360]));

wire [7:0] ens0_layer0_N361_wire = {M0[29], M0[416], M0[562], M0[617], M0[619], M0[631], M0[664], M0[752]};
ens0_layer0_N361 ens0_layer0_N361_inst (.M0(ens0_layer0_N361_wire), .M1(M1[361:361]));

wire [7:0] ens0_layer0_N362_wire = {M0[21], M0[43], M0[477], M0[564], M0[574], M0[586], M0[735], M0[740]};
ens0_layer0_N362 ens0_layer0_N362_inst (.M0(ens0_layer0_N362_wire), .M1(M1[362:362]));

wire [7:0] ens0_layer0_N363_wire = {M0[21], M0[332], M0[396], M0[502], M0[534], M0[623], M0[662], M0[757]};
ens0_layer0_N363 ens0_layer0_N363_inst (.M0(ens0_layer0_N363_wire), .M1(M1[363:363]));

wire [7:0] ens0_layer0_N364_wire = {M0[47], M0[97], M0[316], M0[350], M0[368], M0[389], M0[435], M0[782]};
ens0_layer0_N364 ens0_layer0_N364_inst (.M0(ens0_layer0_N364_wire), .M1(M1[364:364]));

wire [7:0] ens0_layer0_N365_wire = {M0[76], M0[210], M0[250], M0[443], M0[472], M0[539], M0[624], M0[750]};
ens0_layer0_N365 ens0_layer0_N365_inst (.M0(ens0_layer0_N365_wire), .M1(M1[365:365]));

wire [7:0] ens0_layer0_N366_wire = {M0[140], M0[148], M0[289], M0[377], M0[435], M0[506], M0[507], M0[569]};
ens0_layer0_N366 ens0_layer0_N366_inst (.M0(ens0_layer0_N366_wire), .M1(M1[366:366]));

wire [7:0] ens0_layer0_N367_wire = {M0[27], M0[28], M0[247], M0[285], M0[301], M0[316], M0[341], M0[702]};
ens0_layer0_N367 ens0_layer0_N367_inst (.M0(ens0_layer0_N367_wire), .M1(M1[367:367]));

wire [7:0] ens0_layer0_N368_wire = {M0[71], M0[218], M0[235], M0[263], M0[425], M0[585], M0[640], M0[688]};
ens0_layer0_N368 ens0_layer0_N368_inst (.M0(ens0_layer0_N368_wire), .M1(M1[368:368]));

wire [7:0] ens0_layer0_N369_wire = {M0[42], M0[79], M0[86], M0[284], M0[651], M0[679], M0[751], M0[778]};
ens0_layer0_N369 ens0_layer0_N369_inst (.M0(ens0_layer0_N369_wire), .M1(M1[369:369]));

wire [7:0] ens0_layer0_N370_wire = {M0[15], M0[157], M0[258], M0[539], M0[558], M0[583], M0[636], M0[677]};
ens0_layer0_N370 ens0_layer0_N370_inst (.M0(ens0_layer0_N370_wire), .M1(M1[370:370]));

wire [7:0] ens0_layer0_N371_wire = {M0[67], M0[147], M0[151], M0[157], M0[160], M0[336], M0[677], M0[780]};
ens0_layer0_N371 ens0_layer0_N371_inst (.M0(ens0_layer0_N371_wire), .M1(M1[371:371]));

wire [7:0] ens0_layer0_N372_wire = {M0[80], M0[139], M0[272], M0[526], M0[527], M0[659], M0[699], M0[749]};
ens0_layer0_N372 ens0_layer0_N372_inst (.M0(ens0_layer0_N372_wire), .M1(M1[372:372]));

wire [7:0] ens0_layer0_N373_wire = {M0[58], M0[275], M0[438], M0[460], M0[519], M0[559], M0[596], M0[739]};
ens0_layer0_N373 ens0_layer0_N373_inst (.M0(ens0_layer0_N373_wire), .M1(M1[373:373]));

wire [7:0] ens0_layer0_N374_wire = {M0[86], M0[305], M0[327], M0[335], M0[415], M0[520], M0[559], M0[774]};
ens0_layer0_N374 ens0_layer0_N374_inst (.M0(ens0_layer0_N374_wire), .M1(M1[374:374]));

wire [7:0] ens0_layer0_N375_wire = {M0[92], M0[164], M0[177], M0[196], M0[285], M0[414], M0[442], M0[631]};
ens0_layer0_N375 ens0_layer0_N375_inst (.M0(ens0_layer0_N375_wire), .M1(M1[375:375]));

wire [7:0] ens0_layer0_N376_wire = {M0[246], M0[263], M0[330], M0[333], M0[355], M0[470], M0[480], M0[573]};
ens0_layer0_N376 ens0_layer0_N376_inst (.M0(ens0_layer0_N376_wire), .M1(M1[376:376]));

wire [7:0] ens0_layer0_N377_wire = {M0[22], M0[64], M0[247], M0[249], M0[280], M0[294], M0[326], M0[577]};
ens0_layer0_N377 ens0_layer0_N377_inst (.M0(ens0_layer0_N377_wire), .M1(M1[377:377]));

wire [7:0] ens0_layer0_N378_wire = {M0[185], M0[243], M0[328], M0[391], M0[539], M0[557], M0[656], M0[703]};
ens0_layer0_N378 ens0_layer0_N378_inst (.M0(ens0_layer0_N378_wire), .M1(M1[378:378]));

wire [7:0] ens0_layer0_N379_wire = {M0[3], M0[43], M0[516], M0[622], M0[680], M0[690], M0[718], M0[768]};
ens0_layer0_N379 ens0_layer0_N379_inst (.M0(ens0_layer0_N379_wire), .M1(M1[379:379]));

wire [7:0] ens0_layer0_N380_wire = {M0[162], M0[222], M0[456], M0[457], M0[621], M0[656], M0[774], M0[777]};
ens0_layer0_N380 ens0_layer0_N380_inst (.M0(ens0_layer0_N380_wire), .M1(M1[380:380]));

wire [7:0] ens0_layer0_N381_wire = {M0[81], M0[122], M0[274], M0[351], M0[380], M0[385], M0[720], M0[727]};
ens0_layer0_N381 ens0_layer0_N381_inst (.M0(ens0_layer0_N381_wire), .M1(M1[381:381]));

wire [7:0] ens0_layer0_N382_wire = {M0[2], M0[198], M0[200], M0[309], M0[451], M0[482], M0[582], M0[625]};
ens0_layer0_N382 ens0_layer0_N382_inst (.M0(ens0_layer0_N382_wire), .M1(M1[382:382]));

wire [7:0] ens0_layer0_N383_wire = {M0[60], M0[267], M0[284], M0[488], M0[553], M0[597], M0[654], M0[746]};
ens0_layer0_N383 ens0_layer0_N383_inst (.M0(ens0_layer0_N383_wire), .M1(M1[383:383]));

wire [7:0] ens0_layer0_N384_wire = {M0[30], M0[250], M0[501], M0[520], M0[540], M0[561], M0[688], M0[745]};
ens0_layer0_N384 ens0_layer0_N384_inst (.M0(ens0_layer0_N384_wire), .M1(M1[384:384]));

wire [7:0] ens0_layer0_N385_wire = {M0[0], M0[141], M0[148], M0[220], M0[301], M0[331], M0[561], M0[710]};
ens0_layer0_N385 ens0_layer0_N385_inst (.M0(ens0_layer0_N385_wire), .M1(M1[385:385]));

wire [7:0] ens0_layer0_N386_wire = {M0[76], M0[289], M0[570], M0[579], M0[598], M0[653], M0[709], M0[722]};
ens0_layer0_N386 ens0_layer0_N386_inst (.M0(ens0_layer0_N386_wire), .M1(M1[386:386]));

wire [7:0] ens0_layer0_N387_wire = {M0[4], M0[235], M0[309], M0[425], M0[457], M0[593], M0[667], M0[670]};
ens0_layer0_N387 ens0_layer0_N387_inst (.M0(ens0_layer0_N387_wire), .M1(M1[387:387]));

wire [7:0] ens0_layer0_N388_wire = {M0[32], M0[58], M0[84], M0[197], M0[255], M0[299], M0[488], M0[539]};
ens0_layer0_N388 ens0_layer0_N388_inst (.M0(ens0_layer0_N388_wire), .M1(M1[388:388]));

wire [7:0] ens0_layer0_N389_wire = {M0[90], M0[373], M0[393], M0[568], M0[643], M0[665], M0[674], M0[728]};
ens0_layer0_N389 ens0_layer0_N389_inst (.M0(ens0_layer0_N389_wire), .M1(M1[389:389]));

wire [7:0] ens0_layer0_N390_wire = {M0[47], M0[53], M0[94], M0[369], M0[450], M0[594], M0[602], M0[676]};
ens0_layer0_N390 ens0_layer0_N390_inst (.M0(ens0_layer0_N390_wire), .M1(M1[390:390]));

wire [7:0] ens0_layer0_N391_wire = {M0[63], M0[237], M0[296], M0[437], M0[458], M0[546], M0[589], M0[623]};
ens0_layer0_N391 ens0_layer0_N391_inst (.M0(ens0_layer0_N391_wire), .M1(M1[391:391]));

wire [7:0] ens0_layer0_N392_wire = {M0[59], M0[188], M0[210], M0[263], M0[275], M0[448], M0[679], M0[759]};
ens0_layer0_N392 ens0_layer0_N392_inst (.M0(ens0_layer0_N392_wire), .M1(M1[392:392]));

wire [7:0] ens0_layer0_N393_wire = {M0[288], M0[312], M0[324], M0[337], M0[508], M0[510], M0[714], M0[761]};
ens0_layer0_N393 ens0_layer0_N393_inst (.M0(ens0_layer0_N393_wire), .M1(M1[393:393]));

wire [7:0] ens0_layer0_N394_wire = {M0[60], M0[328], M0[516], M0[673], M0[686], M0[747], M0[764], M0[782]};
ens0_layer0_N394 ens0_layer0_N394_inst (.M0(ens0_layer0_N394_wire), .M1(M1[394:394]));

wire [7:0] ens0_layer0_N395_wire = {M0[124], M0[130], M0[366], M0[379], M0[396], M0[443], M0[603], M0[733]};
ens0_layer0_N395 ens0_layer0_N395_inst (.M0(ens0_layer0_N395_wire), .M1(M1[395:395]));

wire [7:0] ens0_layer0_N396_wire = {M0[84], M0[417], M0[504], M0[548], M0[559], M0[592], M0[752], M0[779]};
ens0_layer0_N396 ens0_layer0_N396_inst (.M0(ens0_layer0_N396_wire), .M1(M1[396:396]));

wire [7:0] ens0_layer0_N397_wire = {M0[0], M0[29], M0[119], M0[183], M0[184], M0[409], M0[427], M0[547]};
ens0_layer0_N397 ens0_layer0_N397_inst (.M0(ens0_layer0_N397_wire), .M1(M1[397:397]));

wire [7:0] ens0_layer0_N398_wire = {M0[55], M0[234], M0[272], M0[463], M0[466], M0[488], M0[570], M0[624]};
ens0_layer0_N398 ens0_layer0_N398_inst (.M0(ens0_layer0_N398_wire), .M1(M1[398:398]));

wire [7:0] ens0_layer0_N399_wire = {M0[63], M0[74], M0[123], M0[398], M0[469], M0[529], M0[622], M0[713]};
ens0_layer0_N399 ens0_layer0_N399_inst (.M0(ens0_layer0_N399_wire), .M1(M1[399:399]));

wire [7:0] ens0_layer0_N400_wire = {M0[35], M0[50], M0[71], M0[337], M0[471], M0[497], M0[518], M0[564]};
ens0_layer0_N400 ens0_layer0_N400_inst (.M0(ens0_layer0_N400_wire), .M1(M1[400:400]));

wire [7:0] ens0_layer0_N401_wire = {M0[337], M0[436], M0[438], M0[472], M0[563], M0[664], M0[734], M0[779]};
ens0_layer0_N401 ens0_layer0_N401_inst (.M0(ens0_layer0_N401_wire), .M1(M1[401:401]));

wire [7:0] ens0_layer0_N402_wire = {M0[28], M0[129], M0[155], M0[350], M0[368], M0[425], M0[462], M0[760]};
ens0_layer0_N402 ens0_layer0_N402_inst (.M0(ens0_layer0_N402_wire), .M1(M1[402:402]));

wire [7:0] ens0_layer0_N403_wire = {M0[196], M0[245], M0[263], M0[344], M0[433], M0[463], M0[661], M0[760]};
ens0_layer0_N403 ens0_layer0_N403_inst (.M0(ens0_layer0_N403_wire), .M1(M1[403:403]));

wire [7:0] ens0_layer0_N404_wire = {M0[333], M0[364], M0[398], M0[407], M0[431], M0[515], M0[536], M0[616]};
ens0_layer0_N404 ens0_layer0_N404_inst (.M0(ens0_layer0_N404_wire), .M1(M1[404:404]));

wire [7:0] ens0_layer0_N405_wire = {M0[4], M0[114], M0[126], M0[138], M0[454], M0[504], M0[511], M0[711]};
ens0_layer0_N405 ens0_layer0_N405_inst (.M0(ens0_layer0_N405_wire), .M1(M1[405:405]));

wire [7:0] ens0_layer0_N406_wire = {M0[259], M0[275], M0[308], M0[397], M0[413], M0[500], M0[529], M0[628]};
ens0_layer0_N406 ens0_layer0_N406_inst (.M0(ens0_layer0_N406_wire), .M1(M1[406:406]));

wire [7:0] ens0_layer0_N407_wire = {M0[185], M0[233], M0[246], M0[350], M0[379], M0[486], M0[672], M0[727]};
ens0_layer0_N407 ens0_layer0_N407_inst (.M0(ens0_layer0_N407_wire), .M1(M1[407:407]));

wire [7:0] ens0_layer0_N408_wire = {M0[64], M0[188], M0[336], M0[347], M0[483], M0[590], M0[724], M0[741]};
ens0_layer0_N408 ens0_layer0_N408_inst (.M0(ens0_layer0_N408_wire), .M1(M1[408:408]));

wire [7:0] ens0_layer0_N409_wire = {M0[89], M0[142], M0[155], M0[294], M0[420], M0[473], M0[502], M0[665]};
ens0_layer0_N409 ens0_layer0_N409_inst (.M0(ens0_layer0_N409_wire), .M1(M1[409:409]));

wire [7:0] ens0_layer0_N410_wire = {M0[132], M0[227], M0[257], M0[375], M0[378], M0[414], M0[415], M0[499]};
ens0_layer0_N410 ens0_layer0_N410_inst (.M0(ens0_layer0_N410_wire), .M1(M1[410:410]));

wire [7:0] ens0_layer0_N411_wire = {M0[38], M0[64], M0[86], M0[162], M0[195], M0[215], M0[328], M0[411]};
ens0_layer0_N411 ens0_layer0_N411_inst (.M0(ens0_layer0_N411_wire), .M1(M1[411:411]));

wire [7:0] ens0_layer0_N412_wire = {M0[110], M0[192], M0[318], M0[319], M0[387], M0[467], M0[527], M0[559]};
ens0_layer0_N412 ens0_layer0_N412_inst (.M0(ens0_layer0_N412_wire), .M1(M1[412:412]));

wire [7:0] ens0_layer0_N413_wire = {M0[3], M0[91], M0[128], M0[372], M0[425], M0[513], M0[583], M0[722]};
ens0_layer0_N413 ens0_layer0_N413_inst (.M0(ens0_layer0_N413_wire), .M1(M1[413:413]));

wire [7:0] ens0_layer0_N414_wire = {M0[19], M0[80], M0[117], M0[229], M0[294], M0[299], M0[421], M0[734]};
ens0_layer0_N414 ens0_layer0_N414_inst (.M0(ens0_layer0_N414_wire), .M1(M1[414:414]));

wire [7:0] ens0_layer0_N415_wire = {M0[93], M0[96], M0[265], M0[350], M0[495], M0[543], M0[590], M0[616]};
ens0_layer0_N415 ens0_layer0_N415_inst (.M0(ens0_layer0_N415_wire), .M1(M1[415:415]));

wire [7:0] ens0_layer0_N416_wire = {M0[70], M0[73], M0[237], M0[323], M0[350], M0[401], M0[430], M0[446]};
ens0_layer0_N416 ens0_layer0_N416_inst (.M0(ens0_layer0_N416_wire), .M1(M1[416:416]));

wire [7:0] ens0_layer0_N417_wire = {M0[8], M0[115], M0[133], M0[283], M0[313], M0[370], M0[515], M0[704]};
ens0_layer0_N417 ens0_layer0_N417_inst (.M0(ens0_layer0_N417_wire), .M1(M1[417:417]));

wire [7:0] ens0_layer0_N418_wire = {M0[33], M0[124], M0[138], M0[307], M0[436], M0[479], M0[485], M0[694]};
ens0_layer0_N418 ens0_layer0_N418_inst (.M0(ens0_layer0_N418_wire), .M1(M1[418:418]));

wire [7:0] ens0_layer0_N419_wire = {M0[158], M0[259], M0[335], M0[426], M0[455], M0[488], M0[629], M0[747]};
ens0_layer0_N419 ens0_layer0_N419_inst (.M0(ens0_layer0_N419_wire), .M1(M1[419:419]));

wire [7:0] ens0_layer0_N420_wire = {M0[77], M0[158], M0[248], M0[253], M0[383], M0[595], M0[679], M0[715]};
ens0_layer0_N420 ens0_layer0_N420_inst (.M0(ens0_layer0_N420_wire), .M1(M1[420:420]));

wire [7:0] ens0_layer0_N421_wire = {M0[114], M0[128], M0[339], M0[371], M0[470], M0[553], M0[627], M0[657]};
ens0_layer0_N421 ens0_layer0_N421_inst (.M0(ens0_layer0_N421_wire), .M1(M1[421:421]));

wire [7:0] ens0_layer0_N422_wire = {M0[35], M0[41], M0[396], M0[465], M0[628], M0[716], M0[734], M0[760]};
ens0_layer0_N422 ens0_layer0_N422_inst (.M0(ens0_layer0_N422_wire), .M1(M1[422:422]));

wire [7:0] ens0_layer0_N423_wire = {M0[88], M0[115], M0[262], M0[334], M0[364], M0[458], M0[473], M0[682]};
ens0_layer0_N423 ens0_layer0_N423_inst (.M0(ens0_layer0_N423_wire), .M1(M1[423:423]));

wire [7:0] ens0_layer0_N424_wire = {M0[23], M0[195], M0[224], M0[247], M0[338], M0[417], M0[464], M0[485]};
ens0_layer0_N424 ens0_layer0_N424_inst (.M0(ens0_layer0_N424_wire), .M1(M1[424:424]));

wire [7:0] ens0_layer0_N425_wire = {M0[26], M0[153], M0[370], M0[676], M0[691], M0[698], M0[749], M0[757]};
ens0_layer0_N425 ens0_layer0_N425_inst (.M0(ens0_layer0_N425_wire), .M1(M1[425:425]));

wire [7:0] ens0_layer0_N426_wire = {M0[172], M0[196], M0[201], M0[351], M0[421], M0[435], M0[512], M0[545]};
ens0_layer0_N426 ens0_layer0_N426_inst (.M0(ens0_layer0_N426_wire), .M1(M1[426:426]));

wire [7:0] ens0_layer0_N427_wire = {M0[92], M0[159], M0[330], M0[420], M0[440], M0[496], M0[503], M0[555]};
ens0_layer0_N427 ens0_layer0_N427_inst (.M0(ens0_layer0_N427_wire), .M1(M1[427:427]));

wire [7:0] ens0_layer0_N428_wire = {M0[77], M0[114], M0[139], M0[210], M0[446], M0[487], M0[502], M0[662]};
ens0_layer0_N428 ens0_layer0_N428_inst (.M0(ens0_layer0_N428_wire), .M1(M1[428:428]));

wire [7:0] ens0_layer0_N429_wire = {M0[7], M0[12], M0[240], M0[244], M0[424], M0[435], M0[501], M0[724]};
ens0_layer0_N429 ens0_layer0_N429_inst (.M0(ens0_layer0_N429_wire), .M1(M1[429:429]));

wire [7:0] ens0_layer0_N430_wire = {M0[240], M0[275], M0[328], M0[526], M0[606], M0[609], M0[612], M0[761]};
ens0_layer0_N430 ens0_layer0_N430_inst (.M0(ens0_layer0_N430_wire), .M1(M1[430:430]));

wire [7:0] ens0_layer0_N431_wire = {M0[77], M0[135], M0[234], M0[285], M0[320], M0[568], M0[593], M0[668]};
ens0_layer0_N431 ens0_layer0_N431_inst (.M0(ens0_layer0_N431_wire), .M1(M1[431:431]));

wire [7:0] ens0_layer0_N432_wire = {M0[193], M0[269], M0[277], M0[280], M0[342], M0[569], M0[721], M0[777]};
ens0_layer0_N432 ens0_layer0_N432_inst (.M0(ens0_layer0_N432_wire), .M1(M1[432:432]));

wire [7:0] ens0_layer0_N433_wire = {M0[67], M0[105], M0[296], M0[419], M0[623], M0[626], M0[665], M0[781]};
ens0_layer0_N433 ens0_layer0_N433_inst (.M0(ens0_layer0_N433_wire), .M1(M1[433:433]));

wire [7:0] ens0_layer0_N434_wire = {M0[90], M0[197], M0[230], M0[267], M0[364], M0[593], M0[611], M0[615]};
ens0_layer0_N434 ens0_layer0_N434_inst (.M0(ens0_layer0_N434_wire), .M1(M1[434:434]));

wire [7:0] ens0_layer0_N435_wire = {M0[43], M0[53], M0[353], M0[401], M0[588], M0[617], M0[619], M0[657]};
ens0_layer0_N435 ens0_layer0_N435_inst (.M0(ens0_layer0_N435_wire), .M1(M1[435:435]));

wire [7:0] ens0_layer0_N436_wire = {M0[74], M0[97], M0[147], M0[227], M0[332], M0[584], M0[648], M0[700]};
ens0_layer0_N436 ens0_layer0_N436_inst (.M0(ens0_layer0_N436_wire), .M1(M1[436:436]));

wire [7:0] ens0_layer0_N437_wire = {M0[43], M0[112], M0[154], M0[213], M0[278], M0[377], M0[379], M0[695]};
ens0_layer0_N437 ens0_layer0_N437_inst (.M0(ens0_layer0_N437_wire), .M1(M1[437:437]));

wire [7:0] ens0_layer0_N438_wire = {M0[27], M0[134], M0[179], M0[220], M0[226], M0[428], M0[645], M0[707]};
ens0_layer0_N438 ens0_layer0_N438_inst (.M0(ens0_layer0_N438_wire), .M1(M1[438:438]));

wire [7:0] ens0_layer0_N439_wire = {M0[14], M0[124], M0[282], M0[329], M0[501], M0[521], M0[609], M0[637]};
ens0_layer0_N439 ens0_layer0_N439_inst (.M0(ens0_layer0_N439_wire), .M1(M1[439:439]));

wire [7:0] ens0_layer0_N440_wire = {M0[41], M0[148], M0[165], M0[279], M0[435], M0[462], M0[580], M0[724]};
ens0_layer0_N440 ens0_layer0_N440_inst (.M0(ens0_layer0_N440_wire), .M1(M1[440:440]));

wire [7:0] ens0_layer0_N441_wire = {M0[2], M0[32], M0[345], M0[411], M0[433], M0[438], M0[451], M0[738]};
ens0_layer0_N441 ens0_layer0_N441_inst (.M0(ens0_layer0_N441_wire), .M1(M1[441:441]));

wire [7:0] ens0_layer0_N442_wire = {M0[88], M0[132], M0[227], M0[277], M0[578], M0[670], M0[701], M0[727]};
ens0_layer0_N442 ens0_layer0_N442_inst (.M0(ens0_layer0_N442_wire), .M1(M1[442:442]));

wire [7:0] ens0_layer0_N443_wire = {M0[83], M0[124], M0[240], M0[259], M0[320], M0[378], M0[618], M0[687]};
ens0_layer0_N443 ens0_layer0_N443_inst (.M0(ens0_layer0_N443_wire), .M1(M1[443:443]));

wire [7:0] ens0_layer0_N444_wire = {M0[44], M0[174], M0[243], M0[293], M0[453], M0[469], M0[554], M0[727]};
ens0_layer0_N444 ens0_layer0_N444_inst (.M0(ens0_layer0_N444_wire), .M1(M1[444:444]));

wire [7:0] ens0_layer0_N445_wire = {M0[41], M0[160], M0[246], M0[339], M0[349], M0[423], M0[518], M0[743]};
ens0_layer0_N445 ens0_layer0_N445_inst (.M0(ens0_layer0_N445_wire), .M1(M1[445:445]));

wire [7:0] ens0_layer0_N446_wire = {M0[152], M0[200], M0[202], M0[474], M0[625], M0[633], M0[647], M0[674]};
ens0_layer0_N446 ens0_layer0_N446_inst (.M0(ens0_layer0_N446_wire), .M1(M1[446:446]));

wire [7:0] ens0_layer0_N447_wire = {M0[101], M0[134], M0[205], M0[263], M0[469], M0[477], M0[557], M0[685]};
ens0_layer0_N447 ens0_layer0_N447_inst (.M0(ens0_layer0_N447_wire), .M1(M1[447:447]));

wire [7:0] ens0_layer0_N448_wire = {M0[110], M0[172], M0[221], M0[259], M0[543], M0[652], M0[697], M0[777]};
ens0_layer0_N448 ens0_layer0_N448_inst (.M0(ens0_layer0_N448_wire), .M1(M1[448:448]));

wire [7:0] ens0_layer0_N449_wire = {M0[380], M0[446], M0[510], M0[554], M0[597], M0[682], M0[689], M0[745]};
ens0_layer0_N449 ens0_layer0_N449_inst (.M0(ens0_layer0_N449_wire), .M1(M1[449:449]));

wire [7:0] ens0_layer0_N450_wire = {M0[32], M0[70], M0[91], M0[144], M0[477], M0[546], M0[656], M0[691]};
ens0_layer0_N450 ens0_layer0_N450_inst (.M0(ens0_layer0_N450_wire), .M1(M1[450:450]));

wire [7:0] ens0_layer0_N451_wire = {M0[76], M0[111], M0[168], M0[267], M0[334], M0[388], M0[562], M0[712]};
ens0_layer0_N451 ens0_layer0_N451_inst (.M0(ens0_layer0_N451_wire), .M1(M1[451:451]));

wire [7:0] ens0_layer0_N452_wire = {M0[91], M0[137], M0[142], M0[213], M0[266], M0[336], M0[408], M0[771]};
ens0_layer0_N452 ens0_layer0_N452_inst (.M0(ens0_layer0_N452_wire), .M1(M1[452:452]));

wire [7:0] ens0_layer0_N453_wire = {M0[74], M0[197], M0[253], M0[297], M0[325], M0[333], M0[611], M0[701]};
ens0_layer0_N453 ens0_layer0_N453_inst (.M0(ens0_layer0_N453_wire), .M1(M1[453:453]));

wire [7:0] ens0_layer0_N454_wire = {M0[51], M0[66], M0[123], M0[155], M0[199], M0[430], M0[627], M0[648]};
ens0_layer0_N454 ens0_layer0_N454_inst (.M0(ens0_layer0_N454_wire), .M1(M1[454:454]));

wire [7:0] ens0_layer0_N455_wire = {M0[106], M0[131], M0[285], M0[412], M0[457], M0[595], M0[697], M0[724]};
ens0_layer0_N455 ens0_layer0_N455_inst (.M0(ens0_layer0_N455_wire), .M1(M1[455:455]));

wire [7:0] ens0_layer0_N456_wire = {M0[316], M0[321], M0[351], M0[419], M0[425], M0[436], M0[615], M0[674]};
ens0_layer0_N456 ens0_layer0_N456_inst (.M0(ens0_layer0_N456_wire), .M1(M1[456:456]));

wire [7:0] ens0_layer0_N457_wire = {M0[76], M0[222], M0[295], M0[312], M0[325], M0[334], M0[438], M0[694]};
ens0_layer0_N457 ens0_layer0_N457_inst (.M0(ens0_layer0_N457_wire), .M1(M1[457:457]));

wire [7:0] ens0_layer0_N458_wire = {M0[118], M0[193], M0[318], M0[385], M0[431], M0[563], M0[569], M0[757]};
ens0_layer0_N458 ens0_layer0_N458_inst (.M0(ens0_layer0_N458_wire), .M1(M1[458:458]));

wire [7:0] ens0_layer0_N459_wire = {M0[3], M0[161], M0[414], M0[434], M0[599], M0[621], M0[658], M0[702]};
ens0_layer0_N459 ens0_layer0_N459_inst (.M0(ens0_layer0_N459_wire), .M1(M1[459:459]));

wire [7:0] ens0_layer0_N460_wire = {M0[42], M0[203], M0[279], M0[339], M0[368], M0[445], M0[642], M0[700]};
ens0_layer0_N460 ens0_layer0_N460_inst (.M0(ens0_layer0_N460_wire), .M1(M1[460:460]));

wire [7:0] ens0_layer0_N461_wire = {M0[244], M0[300], M0[333], M0[361], M0[459], M0[544], M0[575], M0[658]};
ens0_layer0_N461 ens0_layer0_N461_inst (.M0(ens0_layer0_N461_wire), .M1(M1[461:461]));

wire [7:0] ens0_layer0_N462_wire = {M0[75], M0[118], M0[352], M0[551], M0[594], M0[623], M0[751], M0[766]};
ens0_layer0_N462 ens0_layer0_N462_inst (.M0(ens0_layer0_N462_wire), .M1(M1[462:462]));

wire [7:0] ens0_layer0_N463_wire = {M0[19], M0[34], M0[93], M0[155], M0[526], M0[541], M0[665], M0[695]};
ens0_layer0_N463 ens0_layer0_N463_inst (.M0(ens0_layer0_N463_wire), .M1(M1[463:463]));

wire [7:0] ens0_layer0_N464_wire = {M0[62], M0[95], M0[165], M0[531], M0[676], M0[704], M0[724], M0[746]};
ens0_layer0_N464 ens0_layer0_N464_inst (.M0(ens0_layer0_N464_wire), .M1(M1[464:464]));

wire [7:0] ens0_layer0_N465_wire = {M0[115], M0[171], M0[212], M0[258], M0[354], M0[381], M0[756], M0[779]};
ens0_layer0_N465 ens0_layer0_N465_inst (.M0(ens0_layer0_N465_wire), .M1(M1[465:465]));

wire [7:0] ens0_layer0_N466_wire = {M0[265], M0[451], M0[455], M0[532], M0[547], M0[576], M0[688], M0[695]};
ens0_layer0_N466 ens0_layer0_N466_inst (.M0(ens0_layer0_N466_wire), .M1(M1[466:466]));

wire [7:0] ens0_layer0_N467_wire = {M0[78], M0[80], M0[106], M0[170], M0[265], M0[352], M0[644], M0[778]};
ens0_layer0_N467 ens0_layer0_N467_inst (.M0(ens0_layer0_N467_wire), .M1(M1[467:467]));

wire [7:0] ens0_layer0_N468_wire = {M0[88], M0[126], M0[201], M0[375], M0[376], M0[544], M0[650], M0[705]};
ens0_layer0_N468 ens0_layer0_N468_inst (.M0(ens0_layer0_N468_wire), .M1(M1[468:468]));

wire [7:0] ens0_layer0_N469_wire = {M0[10], M0[92], M0[154], M0[336], M0[338], M0[569], M0[620], M0[665]};
ens0_layer0_N469 ens0_layer0_N469_inst (.M0(ens0_layer0_N469_wire), .M1(M1[469:469]));

wire [7:0] ens0_layer0_N470_wire = {M0[52], M0[78], M0[138], M0[231], M0[536], M0[543], M0[561], M0[672]};
ens0_layer0_N470 ens0_layer0_N470_inst (.M0(ens0_layer0_N470_wire), .M1(M1[470:470]));

wire [7:0] ens0_layer0_N471_wire = {M0[55], M0[63], M0[130], M0[187], M0[232], M0[252], M0[317], M0[473]};
ens0_layer0_N471 ens0_layer0_N471_inst (.M0(ens0_layer0_N471_wire), .M1(M1[471:471]));

wire [7:0] ens0_layer0_N472_wire = {M0[57], M0[141], M0[168], M0[284], M0[531], M0[608], M0[747], M0[773]};
ens0_layer0_N472 ens0_layer0_N472_inst (.M0(ens0_layer0_N472_wire), .M1(M1[472:472]));

wire [7:0] ens0_layer0_N473_wire = {M0[56], M0[65], M0[151], M0[328], M0[384], M0[397], M0[539], M0[620]};
ens0_layer0_N473 ens0_layer0_N473_inst (.M0(ens0_layer0_N473_wire), .M1(M1[473:473]));

wire [7:0] ens0_layer0_N474_wire = {M0[130], M0[405], M0[530], M0[596], M0[639], M0[704], M0[730], M0[738]};
ens0_layer0_N474 ens0_layer0_N474_inst (.M0(ens0_layer0_N474_wire), .M1(M1[474:474]));

wire [7:0] ens0_layer0_N475_wire = {M0[101], M0[211], M0[303], M0[331], M0[472], M0[556], M0[694], M0[750]};
ens0_layer0_N475 ens0_layer0_N475_inst (.M0(ens0_layer0_N475_wire), .M1(M1[475:475]));

wire [7:0] ens0_layer0_N476_wire = {M0[4], M0[39], M0[63], M0[424], M0[493], M0[515], M0[518], M0[673]};
ens0_layer0_N476 ens0_layer0_N476_inst (.M0(ens0_layer0_N476_wire), .M1(M1[476:476]));

wire [7:0] ens0_layer0_N477_wire = {M0[32], M0[190], M0[250], M0[301], M0[382], M0[483], M0[681], M0[727]};
ens0_layer0_N477 ens0_layer0_N477_inst (.M0(ens0_layer0_N477_wire), .M1(M1[477:477]));

wire [7:0] ens0_layer0_N478_wire = {M0[9], M0[77], M0[225], M0[258], M0[507], M0[512], M0[641], M0[699]};
ens0_layer0_N478 ens0_layer0_N478_inst (.M0(ens0_layer0_N478_wire), .M1(M1[478:478]));

wire [7:0] ens0_layer0_N479_wire = {M0[206], M0[221], M0[342], M0[378], M0[397], M0[609], M0[634], M0[720]};
ens0_layer0_N479 ens0_layer0_N479_inst (.M0(ens0_layer0_N479_wire), .M1(M1[479:479]));

wire [7:0] ens0_layer0_N480_wire = {M0[118], M0[191], M0[219], M0[243], M0[269], M0[682], M0[727], M0[777]};
ens0_layer0_N480 ens0_layer0_N480_inst (.M0(ens0_layer0_N480_wire), .M1(M1[480:480]));

wire [7:0] ens0_layer0_N481_wire = {M0[98], M0[171], M0[240], M0[274], M0[440], M0[614], M0[631], M0[683]};
ens0_layer0_N481 ens0_layer0_N481_inst (.M0(ens0_layer0_N481_wire), .M1(M1[481:481]));

wire [7:0] ens0_layer0_N482_wire = {M0[100], M0[101], M0[176], M0[398], M0[466], M0[560], M0[680], M0[782]};
ens0_layer0_N482 ens0_layer0_N482_inst (.M0(ens0_layer0_N482_wire), .M1(M1[482:482]));

wire [7:0] ens0_layer0_N483_wire = {M0[164], M0[223], M0[224], M0[242], M0[380], M0[571], M0[672], M0[722]};
ens0_layer0_N483 ens0_layer0_N483_inst (.M0(ens0_layer0_N483_wire), .M1(M1[483:483]));

wire [7:0] ens0_layer0_N484_wire = {M0[68], M0[115], M0[165], M0[578], M0[584], M0[626], M0[691], M0[728]};
ens0_layer0_N484 ens0_layer0_N484_inst (.M0(ens0_layer0_N484_wire), .M1(M1[484:484]));

wire [7:0] ens0_layer0_N485_wire = {M0[145], M0[151], M0[187], M0[222], M0[278], M0[347], M0[500], M0[676]};
ens0_layer0_N485 ens0_layer0_N485_inst (.M0(ens0_layer0_N485_wire), .M1(M1[485:485]));

wire [7:0] ens0_layer0_N486_wire = {M0[26], M0[74], M0[163], M0[291], M0[686], M0[688], M0[695], M0[730]};
ens0_layer0_N486 ens0_layer0_N486_inst (.M0(ens0_layer0_N486_wire), .M1(M1[486:486]));

wire [7:0] ens0_layer0_N487_wire = {M0[8], M0[14], M0[182], M0[240], M0[431], M0[473], M0[630], M0[705]};
ens0_layer0_N487 ens0_layer0_N487_inst (.M0(ens0_layer0_N487_wire), .M1(M1[487:487]));

wire [7:0] ens0_layer0_N488_wire = {M0[46], M0[166], M0[366], M0[629], M0[687], M0[719], M0[724], M0[746]};
ens0_layer0_N488 ens0_layer0_N488_inst (.M0(ens0_layer0_N488_wire), .M1(M1[488:488]));

wire [7:0] ens0_layer0_N489_wire = {M0[85], M0[146], M0[151], M0[207], M0[251], M0[312], M0[524], M0[646]};
ens0_layer0_N489 ens0_layer0_N489_inst (.M0(ens0_layer0_N489_wire), .M1(M1[489:489]));

wire [7:0] ens0_layer0_N490_wire = {M0[6], M0[70], M0[120], M0[289], M0[329], M0[332], M0[674], M0[720]};
ens0_layer0_N490 ens0_layer0_N490_inst (.M0(ens0_layer0_N490_wire), .M1(M1[490:490]));

wire [7:0] ens0_layer0_N491_wire = {M0[91], M0[169], M0[209], M0[250], M0[319], M0[421], M0[457], M0[770]};
ens0_layer0_N491 ens0_layer0_N491_inst (.M0(ens0_layer0_N491_wire), .M1(M1[491:491]));

wire [7:0] ens0_layer0_N492_wire = {M0[108], M0[519], M0[534], M0[564], M0[567], M0[594], M0[638], M0[782]};
ens0_layer0_N492 ens0_layer0_N492_inst (.M0(ens0_layer0_N492_wire), .M1(M1[492:492]));

wire [7:0] ens0_layer0_N493_wire = {M0[66], M0[324], M0[371], M0[447], M0[469], M0[528], M0[559], M0[644]};
ens0_layer0_N493 ens0_layer0_N493_inst (.M0(ens0_layer0_N493_wire), .M1(M1[493:493]));

wire [7:0] ens0_layer0_N494_wire = {M0[241], M0[244], M0[372], M0[397], M0[498], M0[529], M0[606], M0[676]};
ens0_layer0_N494 ens0_layer0_N494_inst (.M0(ens0_layer0_N494_wire), .M1(M1[494:494]));

wire [7:0] ens0_layer0_N495_wire = {M0[213], M0[220], M0[256], M0[320], M0[479], M0[525], M0[589], M0[658]};
ens0_layer0_N495 ens0_layer0_N495_inst (.M0(ens0_layer0_N495_wire), .M1(M1[495:495]));

wire [7:0] ens0_layer0_N496_wire = {M0[7], M0[266], M0[335], M0[422], M0[432], M0[500], M0[546], M0[743]};
ens0_layer0_N496 ens0_layer0_N496_inst (.M0(ens0_layer0_N496_wire), .M1(M1[496:496]));

wire [7:0] ens0_layer0_N497_wire = {M0[133], M0[361], M0[379], M0[440], M0[452], M0[635], M0[689], M0[700]};
ens0_layer0_N497 ens0_layer0_N497_inst (.M0(ens0_layer0_N497_wire), .M1(M1[497:497]));

wire [7:0] ens0_layer0_N498_wire = {M0[153], M0[221], M0[272], M0[446], M0[476], M0[593], M0[638], M0[644]};
ens0_layer0_N498 ens0_layer0_N498_inst (.M0(ens0_layer0_N498_wire), .M1(M1[498:498]));

wire [7:0] ens0_layer0_N499_wire = {M0[90], M0[148], M0[249], M0[280], M0[456], M0[634], M0[646], M0[734]};
ens0_layer0_N499 ens0_layer0_N499_inst (.M0(ens0_layer0_N499_wire), .M1(M1[499:499]));

wire [7:0] ens0_layer0_N500_wire = {M0[364], M0[395], M0[445], M0[652], M0[664], M0[698], M0[717], M0[773]};
ens0_layer0_N500 ens0_layer0_N500_inst (.M0(ens0_layer0_N500_wire), .M1(M1[500:500]));

wire [7:0] ens0_layer0_N501_wire = {M0[38], M0[272], M0[362], M0[373], M0[513], M0[613], M0[700], M0[741]};
ens0_layer0_N501 ens0_layer0_N501_inst (.M0(ens0_layer0_N501_wire), .M1(M1[501:501]));

wire [7:0] ens0_layer0_N502_wire = {M0[2], M0[116], M0[118], M0[335], M0[392], M0[484], M0[518], M0[716]};
ens0_layer0_N502 ens0_layer0_N502_inst (.M0(ens0_layer0_N502_wire), .M1(M1[502:502]));

wire [7:0] ens0_layer0_N503_wire = {M0[108], M0[171], M0[337], M0[614], M0[641], M0[715], M0[731], M0[779]};
ens0_layer0_N503 ens0_layer0_N503_inst (.M0(ens0_layer0_N503_wire), .M1(M1[503:503]));

wire [7:0] ens0_layer0_N504_wire = {M0[125], M0[214], M0[268], M0[358], M0[479], M0[713], M0[714], M0[740]};
ens0_layer0_N504 ens0_layer0_N504_inst (.M0(ens0_layer0_N504_wire), .M1(M1[504:504]));

wire [7:0] ens0_layer0_N505_wire = {M0[32], M0[41], M0[53], M0[183], M0[342], M0[506], M0[544], M0[712]};
ens0_layer0_N505 ens0_layer0_N505_inst (.M0(ens0_layer0_N505_wire), .M1(M1[505:505]));

wire [7:0] ens0_layer0_N506_wire = {M0[138], M0[186], M0[206], M0[455], M0[608], M0[674], M0[711], M0[781]};
ens0_layer0_N506 ens0_layer0_N506_inst (.M0(ens0_layer0_N506_wire), .M1(M1[506:506]));

wire [7:0] ens0_layer0_N507_wire = {M0[10], M0[81], M0[94], M0[174], M0[252], M0[256], M0[392], M0[609]};
ens0_layer0_N507 ens0_layer0_N507_inst (.M0(ens0_layer0_N507_wire), .M1(M1[507:507]));

wire [7:0] ens0_layer0_N508_wire = {M0[41], M0[46], M0[371], M0[404], M0[554], M0[566], M0[569], M0[573]};
ens0_layer0_N508 ens0_layer0_N508_inst (.M0(ens0_layer0_N508_wire), .M1(M1[508:508]));

wire [7:0] ens0_layer0_N509_wire = {M0[130], M0[241], M0[251], M0[255], M0[506], M0[585], M0[645], M0[717]};
ens0_layer0_N509 ens0_layer0_N509_inst (.M0(ens0_layer0_N509_wire), .M1(M1[509:509]));

wire [7:0] ens0_layer0_N510_wire = {M0[23], M0[309], M0[367], M0[406], M0[459], M0[560], M0[651], M0[694]};
ens0_layer0_N510 ens0_layer0_N510_inst (.M0(ens0_layer0_N510_wire), .M1(M1[510:510]));

wire [7:0] ens0_layer0_N511_wire = {M0[336], M0[344], M0[387], M0[634], M0[704], M0[724], M0[727], M0[750]};
ens0_layer0_N511 ens0_layer0_N511_inst (.M0(ens0_layer0_N511_wire), .M1(M1[511:511]));

wire [7:0] ens0_layer0_N512_wire = {M0[30], M0[124], M0[165], M0[404], M0[558], M0[567], M0[757], M0[764]};
ens0_layer0_N512 ens0_layer0_N512_inst (.M0(ens0_layer0_N512_wire), .M1(M1[512:512]));

wire [7:0] ens0_layer0_N513_wire = {M0[81], M0[213], M0[263], M0[340], M0[543], M0[627], M0[652], M0[656]};
ens0_layer0_N513 ens0_layer0_N513_inst (.M0(ens0_layer0_N513_wire), .M1(M1[513:513]));

wire [7:0] ens0_layer0_N514_wire = {M0[69], M0[203], M0[285], M0[449], M0[552], M0[660], M0[736], M0[774]};
ens0_layer0_N514 ens0_layer0_N514_inst (.M0(ens0_layer0_N514_wire), .M1(M1[514:514]));

wire [7:0] ens0_layer0_N515_wire = {M0[21], M0[189], M0[293], M0[306], M0[320], M0[445], M0[707], M0[721]};
ens0_layer0_N515 ens0_layer0_N515_inst (.M0(ens0_layer0_N515_wire), .M1(M1[515:515]));

wire [7:0] ens0_layer0_N516_wire = {M0[36], M0[89], M0[192], M0[277], M0[283], M0[503], M0[711], M0[772]};
ens0_layer0_N516 ens0_layer0_N516_inst (.M0(ens0_layer0_N516_wire), .M1(M1[516:516]));

wire [7:0] ens0_layer0_N517_wire = {M0[117], M0[199], M0[204], M0[397], M0[473], M0[684], M0[695], M0[767]};
ens0_layer0_N517 ens0_layer0_N517_inst (.M0(ens0_layer0_N517_wire), .M1(M1[517:517]));

wire [7:0] ens0_layer0_N518_wire = {M0[29], M0[104], M0[135], M0[444], M0[511], M0[599], M0[634], M0[642]};
ens0_layer0_N518 ens0_layer0_N518_inst (.M0(ens0_layer0_N518_wire), .M1(M1[518:518]));

wire [7:0] ens0_layer0_N519_wire = {M0[87], M0[151], M0[247], M0[463], M0[525], M0[661], M0[726], M0[782]};
ens0_layer0_N519 ens0_layer0_N519_inst (.M0(ens0_layer0_N519_wire), .M1(M1[519:519]));

wire [7:0] ens0_layer0_N520_wire = {M0[26], M0[169], M0[249], M0[423], M0[429], M0[477], M0[547], M0[633]};
ens0_layer0_N520 ens0_layer0_N520_inst (.M0(ens0_layer0_N520_wire), .M1(M1[520:520]));

wire [7:0] ens0_layer0_N521_wire = {M0[149], M0[259], M0[371], M0[450], M0[575], M0[624], M0[644], M0[783]};
ens0_layer0_N521 ens0_layer0_N521_inst (.M0(ens0_layer0_N521_wire), .M1(M1[521:521]));

wire [7:0] ens0_layer0_N522_wire = {M0[73], M0[84], M0[101], M0[284], M0[314], M0[430], M0[607], M0[683]};
ens0_layer0_N522 ens0_layer0_N522_inst (.M0(ens0_layer0_N522_wire), .M1(M1[522:522]));

wire [7:0] ens0_layer0_N523_wire = {M0[4], M0[103], M0[238], M0[267], M0[443], M0[454], M0[645], M0[685]};
ens0_layer0_N523 ens0_layer0_N523_inst (.M0(ens0_layer0_N523_wire), .M1(M1[523:523]));

wire [7:0] ens0_layer0_N524_wire = {M0[141], M0[396], M0[420], M0[454], M0[501], M0[563], M0[575], M0[662]};
ens0_layer0_N524 ens0_layer0_N524_inst (.M0(ens0_layer0_N524_wire), .M1(M1[524:524]));

wire [7:0] ens0_layer0_N525_wire = {M0[116], M0[148], M0[162], M0[220], M0[324], M0[534], M0[557], M0[717]};
ens0_layer0_N525 ens0_layer0_N525_inst (.M0(ens0_layer0_N525_wire), .M1(M1[525:525]));

wire [7:0] ens0_layer0_N526_wire = {M0[176], M0[185], M0[210], M0[227], M0[338], M0[344], M0[461], M0[538]};
ens0_layer0_N526 ens0_layer0_N526_inst (.M0(ens0_layer0_N526_wire), .M1(M1[526:526]));

wire [7:0] ens0_layer0_N527_wire = {M0[1], M0[69], M0[138], M0[198], M0[240], M0[269], M0[670], M0[740]};
ens0_layer0_N527 ens0_layer0_N527_inst (.M0(ens0_layer0_N527_wire), .M1(M1[527:527]));

wire [7:0] ens0_layer0_N528_wire = {M0[26], M0[89], M0[104], M0[273], M0[289], M0[516], M0[699], M0[700]};
ens0_layer0_N528 ens0_layer0_N528_inst (.M0(ens0_layer0_N528_wire), .M1(M1[528:528]));

wire [7:0] ens0_layer0_N529_wire = {M0[100], M0[157], M0[158], M0[338], M0[396], M0[588], M0[710], M0[756]};
ens0_layer0_N529 ens0_layer0_N529_inst (.M0(ens0_layer0_N529_wire), .M1(M1[529:529]));

wire [7:0] ens0_layer0_N530_wire = {M0[84], M0[123], M0[126], M0[149], M0[214], M0[454], M0[636], M0[653]};
ens0_layer0_N530 ens0_layer0_N530_inst (.M0(ens0_layer0_N530_wire), .M1(M1[530:530]));

wire [7:0] ens0_layer0_N531_wire = {M0[19], M0[33], M0[228], M0[528], M0[540], M0[605], M0[608], M0[674]};
ens0_layer0_N531 ens0_layer0_N531_inst (.M0(ens0_layer0_N531_wire), .M1(M1[531:531]));

wire [7:0] ens0_layer0_N532_wire = {M0[8], M0[81], M0[125], M0[318], M0[349], M0[518], M0[623], M0[631]};
ens0_layer0_N532 ens0_layer0_N532_inst (.M0(ens0_layer0_N532_wire), .M1(M1[532:532]));

wire [7:0] ens0_layer0_N533_wire = {M0[39], M0[148], M0[166], M0[255], M0[370], M0[394], M0[569], M0[657]};
ens0_layer0_N533 ens0_layer0_N533_inst (.M0(ens0_layer0_N533_wire), .M1(M1[533:533]));

wire [7:0] ens0_layer0_N534_wire = {M0[8], M0[257], M0[440], M0[492], M0[533], M0[686], M0[693], M0[732]};
ens0_layer0_N534 ens0_layer0_N534_inst (.M0(ens0_layer0_N534_wire), .M1(M1[534:534]));

wire [7:0] ens0_layer0_N535_wire = {M0[12], M0[21], M0[72], M0[226], M0[266], M0[430], M0[611], M0[641]};
ens0_layer0_N535 ens0_layer0_N535_inst (.M0(ens0_layer0_N535_wire), .M1(M1[535:535]));

wire [7:0] ens0_layer0_N536_wire = {M0[20], M0[74], M0[129], M0[148], M0[412], M0[447], M0[561], M0[565]};
ens0_layer0_N536 ens0_layer0_N536_inst (.M0(ens0_layer0_N536_wire), .M1(M1[536:536]));

wire [7:0] ens0_layer0_N537_wire = {M0[32], M0[155], M0[165], M0[220], M0[316], M0[369], M0[700], M0[708]};
ens0_layer0_N537 ens0_layer0_N537_inst (.M0(ens0_layer0_N537_wire), .M1(M1[537:537]));

wire [7:0] ens0_layer0_N538_wire = {M0[155], M0[206], M0[330], M0[395], M0[503], M0[581], M0[668], M0[712]};
ens0_layer0_N538 ens0_layer0_N538_inst (.M0(ens0_layer0_N538_wire), .M1(M1[538:538]));

wire [7:0] ens0_layer0_N539_wire = {M0[81], M0[99], M0[328], M0[413], M0[540], M0[544], M0[558], M0[662]};
ens0_layer0_N539 ens0_layer0_N539_inst (.M0(ens0_layer0_N539_wire), .M1(M1[539:539]));

wire [7:0] ens0_layer0_N540_wire = {M0[29], M0[36], M0[216], M0[232], M0[280], M0[428], M0[541], M0[551]};
ens0_layer0_N540 ens0_layer0_N540_inst (.M0(ens0_layer0_N540_wire), .M1(M1[540:540]));

wire [7:0] ens0_layer0_N541_wire = {M0[93], M0[149], M0[214], M0[336], M0[363], M0[380], M0[425], M0[691]};
ens0_layer0_N541 ens0_layer0_N541_inst (.M0(ens0_layer0_N541_wire), .M1(M1[541:541]));

wire [7:0] ens0_layer0_N542_wire = {M0[42], M0[65], M0[262], M0[283], M0[327], M0[359], M0[679], M0[754]};
ens0_layer0_N542 ens0_layer0_N542_inst (.M0(ens0_layer0_N542_wire), .M1(M1[542:542]));

wire [7:0] ens0_layer0_N543_wire = {M0[83], M0[99], M0[150], M0[232], M0[319], M0[464], M0[589], M0[728]};
ens0_layer0_N543 ens0_layer0_N543_inst (.M0(ens0_layer0_N543_wire), .M1(M1[543:543]));

wire [7:0] ens0_layer0_N544_wire = {M0[184], M0[211], M0[221], M0[382], M0[603], M0[628], M0[682], M0[724]};
ens0_layer0_N544 ens0_layer0_N544_inst (.M0(ens0_layer0_N544_wire), .M1(M1[544:544]));

wire [7:0] ens0_layer0_N545_wire = {M0[105], M0[197], M0[229], M0[247], M0[467], M0[534], M0[552], M0[632]};
ens0_layer0_N545 ens0_layer0_N545_inst (.M0(ens0_layer0_N545_wire), .M1(M1[545:545]));

wire [7:0] ens0_layer0_N546_wire = {M0[83], M0[113], M0[262], M0[303], M0[327], M0[428], M0[731], M0[760]};
ens0_layer0_N546 ens0_layer0_N546_inst (.M0(ens0_layer0_N546_wire), .M1(M1[546:546]));

wire [7:0] ens0_layer0_N547_wire = {M0[145], M0[200], M0[291], M0[476], M0[515], M0[536], M0[547], M0[677]};
ens0_layer0_N547 ens0_layer0_N547_inst (.M0(ens0_layer0_N547_wire), .M1(M1[547:547]));

wire [7:0] ens0_layer0_N548_wire = {M0[65], M0[114], M0[127], M0[242], M0[319], M0[599], M0[621], M0[688]};
ens0_layer0_N548 ens0_layer0_N548_inst (.M0(ens0_layer0_N548_wire), .M1(M1[548:548]));

wire [7:0] ens0_layer0_N549_wire = {M0[22], M0[113], M0[115], M0[141], M0[323], M0[714], M0[729], M0[746]};
ens0_layer0_N549 ens0_layer0_N549_inst (.M0(ens0_layer0_N549_wire), .M1(M1[549:549]));

wire [7:0] ens0_layer0_N550_wire = {M0[5], M0[38], M0[75], M0[186], M0[240], M0[417], M0[640], M0[745]};
ens0_layer0_N550 ens0_layer0_N550_inst (.M0(ens0_layer0_N550_wire), .M1(M1[550:550]));

wire [7:0] ens0_layer0_N551_wire = {M0[65], M0[333], M0[342], M0[374], M0[509], M0[627], M0[723], M0[769]};
ens0_layer0_N551 ens0_layer0_N551_inst (.M0(ens0_layer0_N551_wire), .M1(M1[551:551]));

wire [7:0] ens0_layer0_N552_wire = {M0[258], M0[283], M0[335], M0[366], M0[444], M0[499], M0[526], M0[647]};
ens0_layer0_N552 ens0_layer0_N552_inst (.M0(ens0_layer0_N552_wire), .M1(M1[552:552]));

wire [7:0] ens0_layer0_N553_wire = {M0[175], M0[193], M0[234], M0[273], M0[459], M0[522], M0[554], M0[762]};
ens0_layer0_N553 ens0_layer0_N553_inst (.M0(ens0_layer0_N553_wire), .M1(M1[553:553]));

wire [7:0] ens0_layer0_N554_wire = {M0[59], M0[163], M0[300], M0[401], M0[517], M0[573], M0[593], M0[695]};
ens0_layer0_N554 ens0_layer0_N554_inst (.M0(ens0_layer0_N554_wire), .M1(M1[554:554]));

wire [7:0] ens0_layer0_N555_wire = {M0[0], M0[424], M0[469], M0[486], M0[677], M0[685], M0[707], M0[780]};
ens0_layer0_N555 ens0_layer0_N555_inst (.M0(ens0_layer0_N555_wire), .M1(M1[555:555]));

wire [7:0] ens0_layer0_N556_wire = {M0[100], M0[258], M0[315], M0[317], M0[381], M0[429], M0[487], M0[502]};
ens0_layer0_N556 ens0_layer0_N556_inst (.M0(ens0_layer0_N556_wire), .M1(M1[556:556]));

wire [7:0] ens0_layer0_N557_wire = {M0[31], M0[39], M0[158], M0[338], M0[407], M0[434], M0[443], M0[464]};
ens0_layer0_N557 ens0_layer0_N557_inst (.M0(ens0_layer0_N557_wire), .M1(M1[557:557]));

wire [7:0] ens0_layer0_N558_wire = {M0[33], M0[161], M0[169], M0[317], M0[397], M0[459], M0[601], M0[604]};
ens0_layer0_N558 ens0_layer0_N558_inst (.M0(ens0_layer0_N558_wire), .M1(M1[558:558]));

wire [7:0] ens0_layer0_N559_wire = {M0[65], M0[92], M0[149], M0[214], M0[455], M0[553], M0[600], M0[650]};
ens0_layer0_N559 ens0_layer0_N559_inst (.M0(ens0_layer0_N559_wire), .M1(M1[559:559]));

wire [7:0] ens0_layer0_N560_wire = {M0[104], M0[121], M0[157], M0[179], M0[253], M0[330], M0[588], M0[590]};
ens0_layer0_N560 ens0_layer0_N560_inst (.M0(ens0_layer0_N560_wire), .M1(M1[560:560]));

wire [7:0] ens0_layer0_N561_wire = {M0[57], M0[85], M0[254], M0[298], M0[345], M0[367], M0[481], M0[680]};
ens0_layer0_N561 ens0_layer0_N561_inst (.M0(ens0_layer0_N561_wire), .M1(M1[561:561]));

wire [7:0] ens0_layer0_N562_wire = {M0[215], M0[271], M0[285], M0[322], M0[448], M0[588], M0[673], M0[726]};
ens0_layer0_N562 ens0_layer0_N562_inst (.M0(ens0_layer0_N562_wire), .M1(M1[562:562]));

wire [7:0] ens0_layer0_N563_wire = {M0[56], M0[87], M0[365], M0[366], M0[493], M0[672], M0[677], M0[753]};
ens0_layer0_N563 ens0_layer0_N563_inst (.M0(ens0_layer0_N563_wire), .M1(M1[563:563]));

wire [7:0] ens0_layer0_N564_wire = {M0[4], M0[36], M0[310], M0[453], M0[501], M0[666], M0[692], M0[777]};
ens0_layer0_N564 ens0_layer0_N564_inst (.M0(ens0_layer0_N564_wire), .M1(M1[564:564]));

wire [7:0] ens0_layer0_N565_wire = {M0[1], M0[188], M0[252], M0[390], M0[542], M0[604], M0[654], M0[774]};
ens0_layer0_N565 ens0_layer0_N565_inst (.M0(ens0_layer0_N565_wire), .M1(M1[565:565]));

wire [7:0] ens0_layer0_N566_wire = {M0[57], M0[67], M0[195], M0[201], M0[228], M0[470], M0[564], M0[766]};
ens0_layer0_N566 ens0_layer0_N566_inst (.M0(ens0_layer0_N566_wire), .M1(M1[566:566]));

wire [7:0] ens0_layer0_N567_wire = {M0[46], M0[94], M0[106], M0[229], M0[261], M0[277], M0[294], M0[584]};
ens0_layer0_N567 ens0_layer0_N567_inst (.M0(ens0_layer0_N567_wire), .M1(M1[567:567]));

wire [7:0] ens0_layer0_N568_wire = {M0[45], M0[130], M0[131], M0[292], M0[353], M0[464], M0[626], M0[703]};
ens0_layer0_N568 ens0_layer0_N568_inst (.M0(ens0_layer0_N568_wire), .M1(M1[568:568]));

wire [7:0] ens0_layer0_N569_wire = {M0[5], M0[185], M0[316], M0[366], M0[419], M0[583], M0[700], M0[750]};
ens0_layer0_N569 ens0_layer0_N569_inst (.M0(ens0_layer0_N569_wire), .M1(M1[569:569]));

wire [7:0] ens0_layer0_N570_wire = {M0[32], M0[173], M0[212], M0[268], M0[352], M0[385], M0[654], M0[772]};
ens0_layer0_N570 ens0_layer0_N570_inst (.M0(ens0_layer0_N570_wire), .M1(M1[570:570]));

wire [7:0] ens0_layer0_N571_wire = {M0[47], M0[58], M0[180], M0[284], M0[353], M0[407], M0[480], M0[683]};
ens0_layer0_N571 ens0_layer0_N571_inst (.M0(ens0_layer0_N571_wire), .M1(M1[571:571]));

wire [7:0] ens0_layer0_N572_wire = {M0[53], M0[80], M0[301], M0[345], M0[373], M0[535], M0[668], M0[675]};
ens0_layer0_N572 ens0_layer0_N572_inst (.M0(ens0_layer0_N572_wire), .M1(M1[572:572]));

wire [7:0] ens0_layer0_N573_wire = {M0[60], M0[72], M0[259], M0[299], M0[428], M0[460], M0[507], M0[715]};
ens0_layer0_N573 ens0_layer0_N573_inst (.M0(ens0_layer0_N573_wire), .M1(M1[573:573]));

wire [7:0] ens0_layer0_N574_wire = {M0[167], M0[184], M0[247], M0[369], M0[383], M0[388], M0[494], M0[503]};
ens0_layer0_N574 ens0_layer0_N574_inst (.M0(ens0_layer0_N574_wire), .M1(M1[574:574]));

wire [7:0] ens0_layer0_N575_wire = {M0[5], M0[209], M0[294], M0[405], M0[454], M0[519], M0[544], M0[642]};
ens0_layer0_N575 ens0_layer0_N575_inst (.M0(ens0_layer0_N575_wire), .M1(M1[575:575]));

wire [7:0] ens0_layer0_N576_wire = {M0[171], M0[176], M0[213], M0[384], M0[531], M0[648], M0[700], M0[779]};
ens0_layer0_N576 ens0_layer0_N576_inst (.M0(ens0_layer0_N576_wire), .M1(M1[576:576]));

wire [7:0] ens0_layer0_N577_wire = {M0[111], M0[409], M0[442], M0[504], M0[654], M0[664], M0[743], M0[776]};
ens0_layer0_N577 ens0_layer0_N577_inst (.M0(ens0_layer0_N577_wire), .M1(M1[577:577]));

wire [7:0] ens0_layer0_N578_wire = {M0[274], M0[292], M0[320], M0[334], M0[579], M0[597], M0[720], M0[769]};
ens0_layer0_N578 ens0_layer0_N578_inst (.M0(ens0_layer0_N578_wire), .M1(M1[578:578]));

wire [7:0] ens0_layer0_N579_wire = {M0[64], M0[86], M0[106], M0[145], M0[183], M0[238], M0[425], M0[725]};
ens0_layer0_N579 ens0_layer0_N579_inst (.M0(ens0_layer0_N579_wire), .M1(M1[579:579]));

wire [7:0] ens0_layer0_N580_wire = {M0[8], M0[64], M0[103], M0[561], M0[562], M0[631], M0[695], M0[732]};
ens0_layer0_N580 ens0_layer0_N580_inst (.M0(ens0_layer0_N580_wire), .M1(M1[580:580]));

wire [7:0] ens0_layer0_N581_wire = {M0[12], M0[15], M0[116], M0[350], M0[567], M0[613], M0[655], M0[774]};
ens0_layer0_N581 ens0_layer0_N581_inst (.M0(ens0_layer0_N581_wire), .M1(M1[581:581]));

wire [7:0] ens0_layer0_N582_wire = {M0[0], M0[228], M0[460], M0[563], M0[651], M0[724], M0[738], M0[762]};
ens0_layer0_N582 ens0_layer0_N582_inst (.M0(ens0_layer0_N582_wire), .M1(M1[582:582]));

wire [7:0] ens0_layer0_N583_wire = {M0[59], M0[76], M0[78], M0[107], M0[283], M0[561], M0[593], M0[629]};
ens0_layer0_N583 ens0_layer0_N583_inst (.M0(ens0_layer0_N583_wire), .M1(M1[583:583]));

wire [7:0] ens0_layer0_N584_wire = {M0[1], M0[46], M0[103], M0[210], M0[350], M0[483], M0[700], M0[705]};
ens0_layer0_N584 ens0_layer0_N584_inst (.M0(ens0_layer0_N584_wire), .M1(M1[584:584]));

wire [7:0] ens0_layer0_N585_wire = {M0[81], M0[149], M0[283], M0[344], M0[464], M0[626], M0[659], M0[697]};
ens0_layer0_N585 ens0_layer0_N585_inst (.M0(ens0_layer0_N585_wire), .M1(M1[585:585]));

wire [7:0] ens0_layer0_N586_wire = {M0[2], M0[226], M0[230], M0[321], M0[323], M0[348], M0[581], M0[618]};
ens0_layer0_N586 ens0_layer0_N586_inst (.M0(ens0_layer0_N586_wire), .M1(M1[586:586]));

wire [7:0] ens0_layer0_N587_wire = {M0[114], M0[168], M0[181], M0[376], M0[384], M0[481], M0[489], M0[529]};
ens0_layer0_N587 ens0_layer0_N587_inst (.M0(ens0_layer0_N587_wire), .M1(M1[587:587]));

wire [7:0] ens0_layer0_N588_wire = {M0[75], M0[130], M0[219], M0[255], M0[318], M0[352], M0[415], M0[632]};
ens0_layer0_N588 ens0_layer0_N588_inst (.M0(ens0_layer0_N588_wire), .M1(M1[588:588]));

wire [7:0] ens0_layer0_N589_wire = {M0[91], M0[223], M0[473], M0[496], M0[509], M0[645], M0[699], M0[736]};
ens0_layer0_N589 ens0_layer0_N589_inst (.M0(ens0_layer0_N589_wire), .M1(M1[589:589]));

wire [7:0] ens0_layer0_N590_wire = {M0[2], M0[22], M0[263], M0[428], M0[502], M0[545], M0[661], M0[704]};
ens0_layer0_N590 ens0_layer0_N590_inst (.M0(ens0_layer0_N590_wire), .M1(M1[590:590]));

wire [7:0] ens0_layer0_N591_wire = {M0[8], M0[126], M0[273], M0[386], M0[389], M0[550], M0[609], M0[769]};
ens0_layer0_N591 ens0_layer0_N591_inst (.M0(ens0_layer0_N591_wire), .M1(M1[591:591]));

wire [7:0] ens0_layer0_N592_wire = {M0[99], M0[194], M0[296], M0[531], M0[691], M0[701], M0[737], M0[781]};
ens0_layer0_N592 ens0_layer0_N592_inst (.M0(ens0_layer0_N592_wire), .M1(M1[592:592]));

wire [7:0] ens0_layer0_N593_wire = {M0[71], M0[161], M0[192], M0[209], M0[275], M0[319], M0[690], M0[734]};
ens0_layer0_N593 ens0_layer0_N593_inst (.M0(ens0_layer0_N593_wire), .M1(M1[593:593]));

wire [7:0] ens0_layer0_N594_wire = {M0[6], M0[110], M0[129], M0[263], M0[280], M0[403], M0[464], M0[484]};
ens0_layer0_N594 ens0_layer0_N594_inst (.M0(ens0_layer0_N594_wire), .M1(M1[594:594]));

wire [7:0] ens0_layer0_N595_wire = {M0[68], M0[226], M0[369], M0[428], M0[486], M0[509], M0[523], M0[614]};
ens0_layer0_N595 ens0_layer0_N595_inst (.M0(ens0_layer0_N595_wire), .M1(M1[595:595]));

wire [7:0] ens0_layer0_N596_wire = {M0[29], M0[72], M0[75], M0[121], M0[207], M0[384], M0[530], M0[671]};
ens0_layer0_N596 ens0_layer0_N596_inst (.M0(ens0_layer0_N596_wire), .M1(M1[596:596]));

wire [7:0] ens0_layer0_N597_wire = {M0[39], M0[131], M0[215], M0[252], M0[443], M0[514], M0[587], M0[618]};
ens0_layer0_N597 ens0_layer0_N597_inst (.M0(ens0_layer0_N597_wire), .M1(M1[597:597]));

wire [7:0] ens0_layer0_N598_wire = {M0[20], M0[135], M0[358], M0[412], M0[527], M0[582], M0[648], M0[771]};
ens0_layer0_N598 ens0_layer0_N598_inst (.M0(ens0_layer0_N598_wire), .M1(M1[598:598]));

wire [7:0] ens0_layer0_N599_wire = {M0[9], M0[12], M0[151], M0[163], M0[167], M0[353], M0[555], M0[649]};
ens0_layer0_N599 ens0_layer0_N599_inst (.M0(ens0_layer0_N599_wire), .M1(M1[599:599]));

wire [7:0] ens0_layer0_N600_wire = {M0[59], M0[222], M0[269], M0[486], M0[543], M0[629], M0[650], M0[781]};
ens0_layer0_N600 ens0_layer0_N600_inst (.M0(ens0_layer0_N600_wire), .M1(M1[600:600]));

wire [7:0] ens0_layer0_N601_wire = {M0[25], M0[48], M0[71], M0[306], M0[369], M0[511], M0[616], M0[704]};
ens0_layer0_N601 ens0_layer0_N601_inst (.M0(ens0_layer0_N601_wire), .M1(M1[601:601]));

wire [7:0] ens0_layer0_N602_wire = {M0[47], M0[117], M0[188], M0[290], M0[371], M0[430], M0[448], M0[455]};
ens0_layer0_N602 ens0_layer0_N602_inst (.M0(ens0_layer0_N602_wire), .M1(M1[602:602]));

wire [7:0] ens0_layer0_N603_wire = {M0[9], M0[147], M0[186], M0[258], M0[319], M0[361], M0[411], M0[651]};
ens0_layer0_N603 ens0_layer0_N603_inst (.M0(ens0_layer0_N603_wire), .M1(M1[603:603]));

wire [7:0] ens0_layer0_N604_wire = {M0[29], M0[100], M0[114], M0[200], M0[324], M0[387], M0[467], M0[469]};
ens0_layer0_N604 ens0_layer0_N604_inst (.M0(ens0_layer0_N604_wire), .M1(M1[604:604]));

wire [7:0] ens0_layer0_N605_wire = {M0[21], M0[62], M0[83], M0[253], M0[286], M0[573], M0[666], M0[757]};
ens0_layer0_N605 ens0_layer0_N605_inst (.M0(ens0_layer0_N605_wire), .M1(M1[605:605]));

wire [7:0] ens0_layer0_N606_wire = {M0[1], M0[75], M0[137], M0[280], M0[341], M0[379], M0[537], M0[597]};
ens0_layer0_N606 ens0_layer0_N606_inst (.M0(ens0_layer0_N606_wire), .M1(M1[606:606]));

wire [7:0] ens0_layer0_N607_wire = {M0[34], M0[35], M0[104], M0[126], M0[189], M0[545], M0[590], M0[749]};
ens0_layer0_N607 ens0_layer0_N607_inst (.M0(ens0_layer0_N607_wire), .M1(M1[607:607]));

wire [7:0] ens0_layer0_N608_wire = {M0[43], M0[135], M0[196], M0[328], M0[360], M0[412], M0[528], M0[668]};
ens0_layer0_N608 ens0_layer0_N608_inst (.M0(ens0_layer0_N608_wire), .M1(M1[608:608]));

wire [7:0] ens0_layer0_N609_wire = {M0[42], M0[193], M0[235], M0[375], M0[454], M0[490], M0[503], M0[674]};
ens0_layer0_N609 ens0_layer0_N609_inst (.M0(ens0_layer0_N609_wire), .M1(M1[609:609]));

wire [7:0] ens0_layer0_N610_wire = {M0[97], M0[152], M0[155], M0[328], M0[462], M0[520], M0[575], M0[698]};
ens0_layer0_N610 ens0_layer0_N610_inst (.M0(ens0_layer0_N610_wire), .M1(M1[610:610]));

wire [7:0] ens0_layer0_N611_wire = {M0[5], M0[8], M0[33], M0[163], M0[233], M0[373], M0[610], M0[626]};
ens0_layer0_N611 ens0_layer0_N611_inst (.M0(ens0_layer0_N611_wire), .M1(M1[611:611]));

wire [7:0] ens0_layer0_N612_wire = {M0[0], M0[87], M0[129], M0[314], M0[384], M0[538], M0[686], M0[780]};
ens0_layer0_N612 ens0_layer0_N612_inst (.M0(ens0_layer0_N612_wire), .M1(M1[612:612]));

wire [7:0] ens0_layer0_N613_wire = {M0[192], M0[258], M0[365], M0[462], M0[621], M0[695], M0[746], M0[762]};
ens0_layer0_N613 ens0_layer0_N613_inst (.M0(ens0_layer0_N613_wire), .M1(M1[613:613]));

wire [7:0] ens0_layer0_N614_wire = {M0[30], M0[193], M0[249], M0[375], M0[478], M0[480], M0[568], M0[609]};
ens0_layer0_N614 ens0_layer0_N614_inst (.M0(ens0_layer0_N614_wire), .M1(M1[614:614]));

wire [7:0] ens0_layer0_N615_wire = {M0[40], M0[201], M0[223], M0[263], M0[468], M0[486], M0[581], M0[592]};
ens0_layer0_N615 ens0_layer0_N615_inst (.M0(ens0_layer0_N615_wire), .M1(M1[615:615]));

wire [7:0] ens0_layer0_N616_wire = {M0[8], M0[103], M0[118], M0[151], M0[238], M0[401], M0[470], M0[694]};
ens0_layer0_N616 ens0_layer0_N616_inst (.M0(ens0_layer0_N616_wire), .M1(M1[616:616]));

wire [7:0] ens0_layer0_N617_wire = {M0[246], M0[368], M0[441], M0[506], M0[576], M0[702], M0[751], M0[766]};
ens0_layer0_N617 ens0_layer0_N617_inst (.M0(ens0_layer0_N617_wire), .M1(M1[617:617]));

wire [7:0] ens0_layer0_N618_wire = {M0[112], M0[226], M0[242], M0[243], M0[271], M0[348], M0[491], M0[767]};
ens0_layer0_N618 ens0_layer0_N618_inst (.M0(ens0_layer0_N618_wire), .M1(M1[618:618]));

wire [7:0] ens0_layer0_N619_wire = {M0[25], M0[77], M0[214], M0[257], M0[424], M0[479], M0[502], M0[740]};
ens0_layer0_N619 ens0_layer0_N619_inst (.M0(ens0_layer0_N619_wire), .M1(M1[619:619]));

wire [7:0] ens0_layer0_N620_wire = {M0[49], M0[157], M0[162], M0[259], M0[295], M0[400], M0[405], M0[626]};
ens0_layer0_N620 ens0_layer0_N620_inst (.M0(ens0_layer0_N620_wire), .M1(M1[620:620]));

wire [7:0] ens0_layer0_N621_wire = {M0[163], M0[187], M0[254], M0[301], M0[488], M0[494], M0[523], M0[682]};
ens0_layer0_N621 ens0_layer0_N621_inst (.M0(ens0_layer0_N621_wire), .M1(M1[621:621]));

wire [7:0] ens0_layer0_N622_wire = {M0[69], M0[161], M0[181], M0[514], M0[547], M0[551], M0[684], M0[780]};
ens0_layer0_N622 ens0_layer0_N622_inst (.M0(ens0_layer0_N622_wire), .M1(M1[622:622]));

wire [7:0] ens0_layer0_N623_wire = {M0[140], M0[209], M0[264], M0[316], M0[394], M0[464], M0[744], M0[746]};
ens0_layer0_N623 ens0_layer0_N623_inst (.M0(ens0_layer0_N623_wire), .M1(M1[623:623]));

wire [7:0] ens0_layer0_N624_wire = {M0[25], M0[61], M0[143], M0[162], M0[191], M0[438], M0[582], M0[694]};
ens0_layer0_N624 ens0_layer0_N624_inst (.M0(ens0_layer0_N624_wire), .M1(M1[624:624]));

wire [7:0] ens0_layer0_N625_wire = {M0[246], M0[334], M0[483], M0[527], M0[596], M0[660], M0[727], M0[775]};
ens0_layer0_N625 ens0_layer0_N625_inst (.M0(ens0_layer0_N625_wire), .M1(M1[625:625]));

wire [7:0] ens0_layer0_N626_wire = {M0[37], M0[95], M0[100], M0[168], M0[191], M0[284], M0[561], M0[674]};
ens0_layer0_N626 ens0_layer0_N626_inst (.M0(ens0_layer0_N626_wire), .M1(M1[626:626]));

wire [7:0] ens0_layer0_N627_wire = {M0[76], M0[333], M0[497], M0[520], M0[552], M0[637], M0[716], M0[728]};
ens0_layer0_N627 ens0_layer0_N627_inst (.M0(ens0_layer0_N627_wire), .M1(M1[627:627]));

wire [7:0] ens0_layer0_N628_wire = {M0[134], M0[160], M0[202], M0[344], M0[366], M0[495], M0[497], M0[715]};
ens0_layer0_N628 ens0_layer0_N628_inst (.M0(ens0_layer0_N628_wire), .M1(M1[628:628]));

wire [7:0] ens0_layer0_N629_wire = {M0[19], M0[75], M0[107], M0[129], M0[198], M0[442], M0[503], M0[564]};
ens0_layer0_N629 ens0_layer0_N629_inst (.M0(ens0_layer0_N629_wire), .M1(M1[629:629]));

wire [7:0] ens0_layer0_N630_wire = {M0[45], M0[145], M0[291], M0[360], M0[380], M0[597], M0[620], M0[716]};
ens0_layer0_N630 ens0_layer0_N630_inst (.M0(ens0_layer0_N630_wire), .M1(M1[630:630]));

wire [7:0] ens0_layer0_N631_wire = {M0[29], M0[103], M0[120], M0[206], M0[455], M0[523], M0[631], M0[679]};
ens0_layer0_N631 ens0_layer0_N631_inst (.M0(ens0_layer0_N631_wire), .M1(M1[631:631]));

wire [7:0] ens0_layer0_N632_wire = {M0[145], M0[188], M0[461], M0[463], M0[537], M0[541], M0[597], M0[695]};
ens0_layer0_N632 ens0_layer0_N632_inst (.M0(ens0_layer0_N632_wire), .M1(M1[632:632]));

wire [7:0] ens0_layer0_N633_wire = {M0[115], M0[230], M0[342], M0[355], M0[521], M0[530], M0[668], M0[739]};
ens0_layer0_N633 ens0_layer0_N633_inst (.M0(ens0_layer0_N633_wire), .M1(M1[633:633]));

wire [7:0] ens0_layer0_N634_wire = {M0[166], M0[184], M0[221], M0[478], M0[574], M0[614], M0[689], M0[719]};
ens0_layer0_N634 ens0_layer0_N634_inst (.M0(ens0_layer0_N634_wire), .M1(M1[634:634]));

wire [7:0] ens0_layer0_N635_wire = {M0[97], M0[127], M0[136], M0[368], M0[472], M0[474], M0[510], M0[755]};
ens0_layer0_N635 ens0_layer0_N635_inst (.M0(ens0_layer0_N635_wire), .M1(M1[635:635]));

wire [7:0] ens0_layer0_N636_wire = {M0[149], M0[456], M0[458], M0[522], M0[616], M0[631], M0[633], M0[665]};
ens0_layer0_N636 ens0_layer0_N636_inst (.M0(ens0_layer0_N636_wire), .M1(M1[636:636]));

wire [7:0] ens0_layer0_N637_wire = {M0[41], M0[235], M0[281], M0[372], M0[482], M0[534], M0[746], M0[768]};
ens0_layer0_N637 ens0_layer0_N637_inst (.M0(ens0_layer0_N637_wire), .M1(M1[637:637]));

wire [7:0] ens0_layer0_N638_wire = {M0[91], M0[110], M0[291], M0[299], M0[387], M0[443], M0[565], M0[579]};
ens0_layer0_N638 ens0_layer0_N638_inst (.M0(ens0_layer0_N638_wire), .M1(M1[638:638]));

wire [7:0] ens0_layer0_N639_wire = {M0[55], M0[93], M0[106], M0[307], M0[383], M0[511], M0[603], M0[753]};
ens0_layer0_N639 ens0_layer0_N639_inst (.M0(ens0_layer0_N639_wire), .M1(M1[639:639]));

wire [7:0] ens0_layer0_N640_wire = {M0[201], M0[346], M0[350], M0[406], M0[423], M0[441], M0[676], M0[698]};
ens0_layer0_N640 ens0_layer0_N640_inst (.M0(ens0_layer0_N640_wire), .M1(M1[640:640]));

wire [7:0] ens0_layer0_N641_wire = {M0[47], M0[171], M0[177], M0[679], M0[709], M0[771], M0[777], M0[783]};
ens0_layer0_N641 ens0_layer0_N641_inst (.M0(ens0_layer0_N641_wire), .M1(M1[641:641]));

wire [7:0] ens0_layer0_N642_wire = {M0[67], M0[95], M0[100], M0[223], M0[246], M0[324], M0[518], M0[617]};
ens0_layer0_N642 ens0_layer0_N642_inst (.M0(ens0_layer0_N642_wire), .M1(M1[642:642]));

wire [7:0] ens0_layer0_N643_wire = {M0[230], M0[329], M0[430], M0[499], M0[547], M0[576], M0[640], M0[700]};
ens0_layer0_N643 ens0_layer0_N643_inst (.M0(ens0_layer0_N643_wire), .M1(M1[643:643]));

wire [7:0] ens0_layer0_N644_wire = {M0[9], M0[276], M0[347], M0[514], M0[588], M0[617], M0[624], M0[724]};
ens0_layer0_N644 ens0_layer0_N644_inst (.M0(ens0_layer0_N644_wire), .M1(M1[644:644]));

wire [7:0] ens0_layer0_N645_wire = {M0[45], M0[76], M0[264], M0[384], M0[460], M0[502], M0[580], M0[732]};
ens0_layer0_N645 ens0_layer0_N645_inst (.M0(ens0_layer0_N645_wire), .M1(M1[645:645]));

wire [7:0] ens0_layer0_N646_wire = {M0[62], M0[217], M0[238], M0[352], M0[602], M0[642], M0[715], M0[758]};
ens0_layer0_N646 ens0_layer0_N646_inst (.M0(ens0_layer0_N646_wire), .M1(M1[646:646]));

wire [7:0] ens0_layer0_N647_wire = {M0[185], M0[198], M0[374], M0[380], M0[438], M0[586], M0[629], M0[758]};
ens0_layer0_N647 ens0_layer0_N647_inst (.M0(ens0_layer0_N647_wire), .M1(M1[647:647]));

wire [7:0] ens0_layer0_N648_wire = {M0[151], M0[186], M0[281], M0[558], M0[635], M0[640], M0[688], M0[731]};
ens0_layer0_N648 ens0_layer0_N648_inst (.M0(ens0_layer0_N648_wire), .M1(M1[648:648]));

wire [7:0] ens0_layer0_N649_wire = {M0[124], M0[294], M0[348], M0[386], M0[595], M0[699], M0[707], M0[726]};
ens0_layer0_N649 ens0_layer0_N649_inst (.M0(ens0_layer0_N649_wire), .M1(M1[649:649]));

wire [7:0] ens0_layer0_N650_wire = {M0[24], M0[48], M0[100], M0[368], M0[405], M0[429], M0[477], M0[595]};
ens0_layer0_N650 ens0_layer0_N650_inst (.M0(ens0_layer0_N650_wire), .M1(M1[650:650]));

wire [7:0] ens0_layer0_N651_wire = {M0[109], M0[242], M0[348], M0[532], M0[557], M0[580], M0[604], M0[608]};
ens0_layer0_N651 ens0_layer0_N651_inst (.M0(ens0_layer0_N651_wire), .M1(M1[651:651]));

wire [7:0] ens0_layer0_N652_wire = {M0[16], M0[117], M0[236], M0[518], M0[736], M0[770], M0[782], M0[783]};
ens0_layer0_N652 ens0_layer0_N652_inst (.M0(ens0_layer0_N652_wire), .M1(M1[652:652]));

wire [7:0] ens0_layer0_N653_wire = {M0[28], M0[50], M0[126], M0[187], M0[239], M0[595], M0[626], M0[781]};
ens0_layer0_N653 ens0_layer0_N653_inst (.M0(ens0_layer0_N653_wire), .M1(M1[653:653]));

wire [7:0] ens0_layer0_N654_wire = {M0[90], M0[167], M0[207], M0[314], M0[345], M0[430], M0[486], M0[589]};
ens0_layer0_N654 ens0_layer0_N654_inst (.M0(ens0_layer0_N654_wire), .M1(M1[654:654]));

wire [7:0] ens0_layer0_N655_wire = {M0[105], M0[188], M0[230], M0[317], M0[465], M0[513], M0[676], M0[712]};
ens0_layer0_N655 ens0_layer0_N655_inst (.M0(ens0_layer0_N655_wire), .M1(M1[655:655]));

wire [7:0] ens0_layer0_N656_wire = {M0[284], M0[290], M0[295], M0[310], M0[400], M0[432], M0[437], M0[719]};
ens0_layer0_N656 ens0_layer0_N656_inst (.M0(ens0_layer0_N656_wire), .M1(M1[656:656]));

wire [7:0] ens0_layer0_N657_wire = {M0[156], M0[165], M0[263], M0[319], M0[385], M0[485], M0[562], M0[721]};
ens0_layer0_N657 ens0_layer0_N657_inst (.M0(ens0_layer0_N657_wire), .M1(M1[657:657]));

wire [7:0] ens0_layer0_N658_wire = {M0[9], M0[48], M0[206], M0[360], M0[700], M0[739], M0[755], M0[765]};
ens0_layer0_N658 ens0_layer0_N658_inst (.M0(ens0_layer0_N658_wire), .M1(M1[658:658]));

wire [7:0] ens0_layer0_N659_wire = {M0[269], M0[320], M0[401], M0[472], M0[575], M0[678], M0[681], M0[776]};
ens0_layer0_N659 ens0_layer0_N659_inst (.M0(ens0_layer0_N659_wire), .M1(M1[659:659]));

wire [7:0] ens0_layer0_N660_wire = {M0[59], M0[201], M0[208], M0[213], M0[389], M0[476], M0[677], M0[682]};
ens0_layer0_N660 ens0_layer0_N660_inst (.M0(ens0_layer0_N660_wire), .M1(M1[660:660]));

wire [7:0] ens0_layer0_N661_wire = {M0[87], M0[134], M0[274], M0[317], M0[394], M0[400], M0[418], M0[728]};
ens0_layer0_N661 ens0_layer0_N661_inst (.M0(ens0_layer0_N661_wire), .M1(M1[661:661]));

wire [7:0] ens0_layer0_N662_wire = {M0[28], M0[40], M0[143], M0[223], M0[437], M0[568], M0[573], M0[736]};
ens0_layer0_N662 ens0_layer0_N662_inst (.M0(ens0_layer0_N662_wire), .M1(M1[662:662]));

wire [7:0] ens0_layer0_N663_wire = {M0[135], M0[193], M0[352], M0[377], M0[447], M0[548], M0[612], M0[631]};
ens0_layer0_N663 ens0_layer0_N663_inst (.M0(ens0_layer0_N663_wire), .M1(M1[663:663]));

wire [7:0] ens0_layer0_N664_wire = {M0[34], M0[41], M0[81], M0[115], M0[228], M0[336], M0[581], M0[709]};
ens0_layer0_N664 ens0_layer0_N664_inst (.M0(ens0_layer0_N664_wire), .M1(M1[664:664]));

wire [7:0] ens0_layer0_N665_wire = {M0[183], M0[203], M0[246], M0[279], M0[323], M0[384], M0[466], M0[713]};
ens0_layer0_N665 ens0_layer0_N665_inst (.M0(ens0_layer0_N665_wire), .M1(M1[665:665]));

wire [7:0] ens0_layer0_N666_wire = {M0[112], M0[128], M0[399], M0[472], M0[481], M0[511], M0[513], M0[575]};
ens0_layer0_N666 ens0_layer0_N666_inst (.M0(ens0_layer0_N666_wire), .M1(M1[666:666]));

wire [7:0] ens0_layer0_N667_wire = {M0[99], M0[165], M0[247], M0[302], M0[331], M0[447], M0[581], M0[617]};
ens0_layer0_N667 ens0_layer0_N667_inst (.M0(ens0_layer0_N667_wire), .M1(M1[667:667]));

wire [7:0] ens0_layer0_N668_wire = {M0[275], M0[435], M0[580], M0[616], M0[678], M0[696], M0[733], M0[734]};
ens0_layer0_N668 ens0_layer0_N668_inst (.M0(ens0_layer0_N668_wire), .M1(M1[668:668]));

wire [7:0] ens0_layer0_N669_wire = {M0[99], M0[220], M0[290], M0[322], M0[485], M0[628], M0[717], M0[776]};
ens0_layer0_N669 ens0_layer0_N669_inst (.M0(ens0_layer0_N669_wire), .M1(M1[669:669]));

wire [7:0] ens0_layer0_N670_wire = {M0[169], M0[276], M0[395], M0[526], M0[588], M0[608], M0[652], M0[718]};
ens0_layer0_N670 ens0_layer0_N670_inst (.M0(ens0_layer0_N670_wire), .M1(M1[670:670]));

wire [7:0] ens0_layer0_N671_wire = {M0[55], M0[207], M0[324], M0[510], M0[574], M0[617], M0[646], M0[699]};
ens0_layer0_N671 ens0_layer0_N671_inst (.M0(ens0_layer0_N671_wire), .M1(M1[671:671]));

wire [7:0] ens0_layer0_N672_wire = {M0[80], M0[87], M0[96], M0[507], M0[644], M0[668], M0[687], M0[744]};
ens0_layer0_N672 ens0_layer0_N672_inst (.M0(ens0_layer0_N672_wire), .M1(M1[672:672]));

wire [7:0] ens0_layer0_N673_wire = {M0[12], M0[124], M0[199], M0[216], M0[403], M0[552], M0[613], M0[782]};
ens0_layer0_N673 ens0_layer0_N673_inst (.M0(ens0_layer0_N673_wire), .M1(M1[673:673]));

wire [7:0] ens0_layer0_N674_wire = {M0[260], M0[332], M0[393], M0[404], M0[492], M0[569], M0[620], M0[698]};
ens0_layer0_N674 ens0_layer0_N674_inst (.M0(ens0_layer0_N674_wire), .M1(M1[674:674]));

wire [7:0] ens0_layer0_N675_wire = {M0[6], M0[211], M0[471], M0[515], M0[602], M0[631], M0[654], M0[753]};
ens0_layer0_N675 ens0_layer0_N675_inst (.M0(ens0_layer0_N675_wire), .M1(M1[675:675]));

wire [7:0] ens0_layer0_N676_wire = {M0[120], M0[220], M0[435], M0[555], M0[574], M0[609], M0[625], M0[737]};
ens0_layer0_N676 ens0_layer0_N676_inst (.M0(ens0_layer0_N676_wire), .M1(M1[676:676]));

wire [7:0] ens0_layer0_N677_wire = {M0[15], M0[145], M0[259], M0[364], M0[491], M0[494], M0[523], M0[548]};
ens0_layer0_N677 ens0_layer0_N677_inst (.M0(ens0_layer0_N677_wire), .M1(M1[677:677]));

wire [7:0] ens0_layer0_N678_wire = {M0[34], M0[373], M0[431], M0[436], M0[568], M0[711], M0[714], M0[782]};
ens0_layer0_N678 ens0_layer0_N678_inst (.M0(ens0_layer0_N678_wire), .M1(M1[678:678]));

wire [7:0] ens0_layer0_N679_wire = {M0[135], M0[199], M0[331], M0[346], M0[621], M0[652], M0[690], M0[705]};
ens0_layer0_N679 ens0_layer0_N679_inst (.M0(ens0_layer0_N679_wire), .M1(M1[679:679]));

wire [7:0] ens0_layer0_N680_wire = {M0[6], M0[47], M0[166], M0[270], M0[304], M0[497], M0[508], M0[641]};
ens0_layer0_N680 ens0_layer0_N680_inst (.M0(ens0_layer0_N680_wire), .M1(M1[680:680]));

wire [7:0] ens0_layer0_N681_wire = {M0[248], M0[341], M0[482], M0[526], M0[557], M0[632], M0[634], M0[756]};
ens0_layer0_N681 ens0_layer0_N681_inst (.M0(ens0_layer0_N681_wire), .M1(M1[681:681]));

wire [7:0] ens0_layer0_N682_wire = {M0[125], M0[184], M0[236], M0[258], M0[472], M0[501], M0[592], M0[718]};
ens0_layer0_N682 ens0_layer0_N682_inst (.M0(ens0_layer0_N682_wire), .M1(M1[682:682]));

wire [7:0] ens0_layer0_N683_wire = {M0[43], M0[383], M0[417], M0[477], M0[545], M0[605], M0[613], M0[778]};
ens0_layer0_N683 ens0_layer0_N683_inst (.M0(ens0_layer0_N683_wire), .M1(M1[683:683]));

wire [7:0] ens0_layer0_N684_wire = {M0[28], M0[174], M0[344], M0[353], M0[365], M0[558], M0[589], M0[733]};
ens0_layer0_N684 ens0_layer0_N684_inst (.M0(ens0_layer0_N684_wire), .M1(M1[684:684]));

wire [7:0] ens0_layer0_N685_wire = {M0[18], M0[81], M0[155], M0[476], M0[521], M0[628], M0[646], M0[781]};
ens0_layer0_N685 ens0_layer0_N685_inst (.M0(ens0_layer0_N685_wire), .M1(M1[685:685]));

wire [7:0] ens0_layer0_N686_wire = {M0[83], M0[128], M0[142], M0[147], M0[478], M0[487], M0[685], M0[706]};
ens0_layer0_N686 ens0_layer0_N686_inst (.M0(ens0_layer0_N686_wire), .M1(M1[686:686]));

wire [7:0] ens0_layer0_N687_wire = {M0[36], M0[102], M0[380], M0[457], M0[465], M0[548], M0[560], M0[575]};
ens0_layer0_N687 ens0_layer0_N687_inst (.M0(ens0_layer0_N687_wire), .M1(M1[687:687]));

wire [7:0] ens0_layer0_N688_wire = {M0[2], M0[107], M0[334], M0[596], M0[608], M0[619], M0[686], M0[744]};
ens0_layer0_N688 ens0_layer0_N688_inst (.M0(ens0_layer0_N688_wire), .M1(M1[688:688]));

wire [7:0] ens0_layer0_N689_wire = {M0[24], M0[45], M0[77], M0[312], M0[379], M0[495], M0[725], M0[773]};
ens0_layer0_N689 ens0_layer0_N689_inst (.M0(ens0_layer0_N689_wire), .M1(M1[689:689]));

wire [7:0] ens0_layer0_N690_wire = {M0[13], M0[119], M0[314], M0[371], M0[462], M0[492], M0[501], M0[758]};
ens0_layer0_N690 ens0_layer0_N690_inst (.M0(ens0_layer0_N690_wire), .M1(M1[690:690]));

wire [7:0] ens0_layer0_N691_wire = {M0[20], M0[28], M0[37], M0[79], M0[114], M0[192], M0[337], M0[395]};
ens0_layer0_N691 ens0_layer0_N691_inst (.M0(ens0_layer0_N691_wire), .M1(M1[691:691]));

wire [7:0] ens0_layer0_N692_wire = {M0[11], M0[73], M0[151], M0[160], M0[246], M0[274], M0[559], M0[590]};
ens0_layer0_N692 ens0_layer0_N692_inst (.M0(ens0_layer0_N692_wire), .M1(M1[692:692]));

wire [7:0] ens0_layer0_N693_wire = {M0[15], M0[17], M0[31], M0[151], M0[301], M0[319], M0[672], M0[698]};
ens0_layer0_N693 ens0_layer0_N693_inst (.M0(ens0_layer0_N693_wire), .M1(M1[693:693]));

wire [7:0] ens0_layer0_N694_wire = {M0[63], M0[171], M0[207], M0[569], M0[580], M0[589], M0[672], M0[732]};
ens0_layer0_N694 ens0_layer0_N694_inst (.M0(ens0_layer0_N694_wire), .M1(M1[694:694]));

wire [7:0] ens0_layer0_N695_wire = {M0[0], M0[149], M0[191], M0[208], M0[433], M0[636], M0[638], M0[756]};
ens0_layer0_N695 ens0_layer0_N695_inst (.M0(ens0_layer0_N695_wire), .M1(M1[695:695]));

wire [7:0] ens0_layer0_N696_wire = {M0[229], M0[286], M0[337], M0[407], M0[423], M0[619], M0[649], M0[778]};
ens0_layer0_N696 ens0_layer0_N696_inst (.M0(ens0_layer0_N696_wire), .M1(M1[696:696]));

wire [7:0] ens0_layer0_N697_wire = {M0[176], M0[180], M0[494], M0[506], M0[654], M0[732], M0[739], M0[740]};
ens0_layer0_N697 ens0_layer0_N697_inst (.M0(ens0_layer0_N697_wire), .M1(M1[697:697]));

wire [7:0] ens0_layer0_N698_wire = {M0[162], M0[254], M0[276], M0[294], M0[410], M0[425], M0[509], M0[552]};
ens0_layer0_N698 ens0_layer0_N698_inst (.M0(ens0_layer0_N698_wire), .M1(M1[698:698]));

wire [7:0] ens0_layer0_N699_wire = {M0[45], M0[129], M0[231], M0[281], M0[429], M0[511], M0[637], M0[728]};
ens0_layer0_N699 ens0_layer0_N699_inst (.M0(ens0_layer0_N699_wire), .M1(M1[699:699]));

wire [7:0] ens0_layer0_N700_wire = {M0[62], M0[112], M0[254], M0[278], M0[456], M0[465], M0[652], M0[744]};
ens0_layer0_N700 ens0_layer0_N700_inst (.M0(ens0_layer0_N700_wire), .M1(M1[700:700]));

wire [7:0] ens0_layer0_N701_wire = {M0[61], M0[177], M0[246], M0[403], M0[456], M0[489], M0[591], M0[707]};
ens0_layer0_N701 ens0_layer0_N701_inst (.M0(ens0_layer0_N701_wire), .M1(M1[701:701]));

wire [7:0] ens0_layer0_N702_wire = {M0[51], M0[77], M0[83], M0[199], M0[205], M0[363], M0[448], M0[628]};
ens0_layer0_N702 ens0_layer0_N702_inst (.M0(ens0_layer0_N702_wire), .M1(M1[702:702]));

wire [7:0] ens0_layer0_N703_wire = {M0[23], M0[40], M0[258], M0[397], M0[506], M0[565], M0[676], M0[726]};
ens0_layer0_N703 ens0_layer0_N703_inst (.M0(ens0_layer0_N703_wire), .M1(M1[703:703]));

wire [7:0] ens0_layer0_N704_wire = {M0[92], M0[503], M0[511], M0[528], M0[552], M0[560], M0[624], M0[719]};
ens0_layer0_N704 ens0_layer0_N704_inst (.M0(ens0_layer0_N704_wire), .M1(M1[704:704]));

wire [7:0] ens0_layer0_N705_wire = {M0[10], M0[35], M0[262], M0[305], M0[311], M0[368], M0[438], M0[780]};
ens0_layer0_N705 ens0_layer0_N705_inst (.M0(ens0_layer0_N705_wire), .M1(M1[705:705]));

wire [7:0] ens0_layer0_N706_wire = {M0[81], M0[100], M0[146], M0[255], M0[430], M0[610], M0[649], M0[656]};
ens0_layer0_N706 ens0_layer0_N706_inst (.M0(ens0_layer0_N706_wire), .M1(M1[706:706]));

wire [7:0] ens0_layer0_N707_wire = {M0[12], M0[45], M0[193], M0[202], M0[208], M0[249], M0[343], M0[672]};
ens0_layer0_N707 ens0_layer0_N707_inst (.M0(ens0_layer0_N707_wire), .M1(M1[707:707]));

wire [7:0] ens0_layer0_N708_wire = {M0[106], M0[144], M0[236], M0[459], M0[493], M0[533], M0[543], M0[702]};
ens0_layer0_N708 ens0_layer0_N708_inst (.M0(ens0_layer0_N708_wire), .M1(M1[708:708]));

wire [7:0] ens0_layer0_N709_wire = {M0[60], M0[110], M0[225], M0[271], M0[292], M0[475], M0[552], M0[591]};
ens0_layer0_N709 ens0_layer0_N709_inst (.M0(ens0_layer0_N709_wire), .M1(M1[709:709]));

wire [7:0] ens0_layer0_N710_wire = {M0[87], M0[122], M0[147], M0[180], M0[202], M0[427], M0[432], M0[743]};
ens0_layer0_N710 ens0_layer0_N710_inst (.M0(ens0_layer0_N710_wire), .M1(M1[710:710]));

wire [7:0] ens0_layer0_N711_wire = {M0[34], M0[168], M0[186], M0[202], M0[338], M0[357], M0[595], M0[744]};
ens0_layer0_N711 ens0_layer0_N711_inst (.M0(ens0_layer0_N711_wire), .M1(M1[711:711]));

wire [7:0] ens0_layer0_N712_wire = {M0[83], M0[150], M0[317], M0[350], M0[418], M0[512], M0[590], M0[724]};
ens0_layer0_N712 ens0_layer0_N712_inst (.M0(ens0_layer0_N712_wire), .M1(M1[712:712]));

wire [7:0] ens0_layer0_N713_wire = {M0[7], M0[8], M0[56], M0[63], M0[581], M0[604], M0[641], M0[741]};
ens0_layer0_N713 ens0_layer0_N713_inst (.M0(ens0_layer0_N713_wire), .M1(M1[713:713]));

wire [7:0] ens0_layer0_N714_wire = {M0[17], M0[62], M0[83], M0[206], M0[302], M0[364], M0[586], M0[783]};
ens0_layer0_N714 ens0_layer0_N714_inst (.M0(ens0_layer0_N714_wire), .M1(M1[714:714]));

wire [7:0] ens0_layer0_N715_wire = {M0[41], M0[270], M0[324], M0[386], M0[429], M0[466], M0[518], M0[526]};
ens0_layer0_N715 ens0_layer0_N715_inst (.M0(ens0_layer0_N715_wire), .M1(M1[715:715]));

wire [7:0] ens0_layer0_N716_wire = {M0[216], M0[253], M0[364], M0[380], M0[668], M0[672], M0[676], M0[684]};
ens0_layer0_N716 ens0_layer0_N716_inst (.M0(ens0_layer0_N716_wire), .M1(M1[716:716]));

wire [7:0] ens0_layer0_N717_wire = {M0[22], M0[44], M0[104], M0[233], M0[291], M0[491], M0[543], M0[772]};
ens0_layer0_N717 ens0_layer0_N717_inst (.M0(ens0_layer0_N717_wire), .M1(M1[717:717]));

wire [7:0] ens0_layer0_N718_wire = {M0[124], M0[247], M0[296], M0[297], M0[321], M0[371], M0[557], M0[588]};
ens0_layer0_N718 ens0_layer0_N718_inst (.M0(ens0_layer0_N718_wire), .M1(M1[718:718]));

wire [7:0] ens0_layer0_N719_wire = {M0[34], M0[44], M0[169], M0[235], M0[243], M0[267], M0[448], M0[635]};
ens0_layer0_N719 ens0_layer0_N719_inst (.M0(ens0_layer0_N719_wire), .M1(M1[719:719]));

wire [7:0] ens0_layer0_N720_wire = {M0[60], M0[165], M0[362], M0[488], M0[512], M0[519], M0[521], M0[534]};
ens0_layer0_N720 ens0_layer0_N720_inst (.M0(ens0_layer0_N720_wire), .M1(M1[720:720]));

wire [7:0] ens0_layer0_N721_wire = {M0[294], M0[330], M0[344], M0[363], M0[369], M0[430], M0[713], M0[742]};
ens0_layer0_N721 ens0_layer0_N721_inst (.M0(ens0_layer0_N721_wire), .M1(M1[721:721]));

wire [7:0] ens0_layer0_N722_wire = {M0[1], M0[58], M0[91], M0[138], M0[223], M0[529], M0[648], M0[702]};
ens0_layer0_N722 ens0_layer0_N722_inst (.M0(ens0_layer0_N722_wire), .M1(M1[722:722]));

wire [7:0] ens0_layer0_N723_wire = {M0[89], M0[314], M0[438], M0[471], M0[480], M0[509], M0[568], M0[705]};
ens0_layer0_N723 ens0_layer0_N723_inst (.M0(ens0_layer0_N723_wire), .M1(M1[723:723]));

wire [7:0] ens0_layer0_N724_wire = {M0[96], M0[174], M0[262], M0[309], M0[389], M0[523], M0[528], M0[710]};
ens0_layer0_N724 ens0_layer0_N724_inst (.M0(ens0_layer0_N724_wire), .M1(M1[724:724]));

wire [7:0] ens0_layer0_N725_wire = {M0[48], M0[110], M0[230], M0[324], M0[377], M0[430], M0[445], M0[612]};
ens0_layer0_N725 ens0_layer0_N725_inst (.M0(ens0_layer0_N725_wire), .M1(M1[725:725]));

wire [7:0] ens0_layer0_N726_wire = {M0[148], M0[297], M0[329], M0[471], M0[486], M0[564], M0[570], M0[722]};
ens0_layer0_N726 ens0_layer0_N726_inst (.M0(ens0_layer0_N726_wire), .M1(M1[726:726]));

wire [7:0] ens0_layer0_N727_wire = {M0[37], M0[96], M0[140], M0[173], M0[377], M0[402], M0[447], M0[461]};
ens0_layer0_N727 ens0_layer0_N727_inst (.M0(ens0_layer0_N727_wire), .M1(M1[727:727]));

wire [7:0] ens0_layer0_N728_wire = {M0[242], M0[299], M0[359], M0[387], M0[392], M0[460], M0[493], M0[715]};
ens0_layer0_N728 ens0_layer0_N728_inst (.M0(ens0_layer0_N728_wire), .M1(M1[728:728]));

wire [7:0] ens0_layer0_N729_wire = {M0[15], M0[118], M0[210], M0[281], M0[466], M0[527], M0[537], M0[743]};
ens0_layer0_N729 ens0_layer0_N729_inst (.M0(ens0_layer0_N729_wire), .M1(M1[729:729]));

wire [7:0] ens0_layer0_N730_wire = {M0[190], M0[333], M0[337], M0[437], M0[442], M0[667], M0[695], M0[779]};
ens0_layer0_N730 ens0_layer0_N730_inst (.M0(ens0_layer0_N730_wire), .M1(M1[730:730]));

wire [7:0] ens0_layer0_N731_wire = {M0[113], M0[150], M0[418], M0[452], M0[474], M0[561], M0[587], M0[724]};
ens0_layer0_N731 ens0_layer0_N731_inst (.M0(ens0_layer0_N731_wire), .M1(M1[731:731]));

wire [7:0] ens0_layer0_N732_wire = {M0[47], M0[53], M0[117], M0[151], M0[181], M0[255], M0[354], M0[659]};
ens0_layer0_N732 ens0_layer0_N732_inst (.M0(ens0_layer0_N732_wire), .M1(M1[732:732]));

wire [7:0] ens0_layer0_N733_wire = {M0[36], M0[202], M0[249], M0[534], M0[556], M0[683], M0[773], M0[774]};
ens0_layer0_N733 ens0_layer0_N733_inst (.M0(ens0_layer0_N733_wire), .M1(M1[733:733]));

wire [7:0] ens0_layer0_N734_wire = {M0[222], M0[299], M0[489], M0[508], M0[522], M0[535], M0[726], M0[764]};
ens0_layer0_N734 ens0_layer0_N734_inst (.M0(ens0_layer0_N734_wire), .M1(M1[734:734]));

wire [7:0] ens0_layer0_N735_wire = {M0[49], M0[342], M0[427], M0[664], M0[697], M0[700], M0[759], M0[766]};
ens0_layer0_N735 ens0_layer0_N735_inst (.M0(ens0_layer0_N735_wire), .M1(M1[735:735]));

wire [7:0] ens0_layer0_N736_wire = {M0[72], M0[100], M0[140], M0[269], M0[301], M0[486], M0[541], M0[768]};
ens0_layer0_N736 ens0_layer0_N736_inst (.M0(ens0_layer0_N736_wire), .M1(M1[736:736]));

wire [7:0] ens0_layer0_N737_wire = {M0[3], M0[37], M0[144], M0[162], M0[203], M0[309], M0[512], M0[779]};
ens0_layer0_N737 ens0_layer0_N737_inst (.M0(ens0_layer0_N737_wire), .M1(M1[737:737]));

wire [7:0] ens0_layer0_N738_wire = {M0[138], M0[175], M0[316], M0[335], M0[468], M0[525], M0[580], M0[616]};
ens0_layer0_N738 ens0_layer0_N738_inst (.M0(ens0_layer0_N738_wire), .M1(M1[738:738]));

wire [7:0] ens0_layer0_N739_wire = {M0[41], M0[54], M0[197], M0[211], M0[320], M0[616], M0[723], M0[732]};
ens0_layer0_N739 ens0_layer0_N739_inst (.M0(ens0_layer0_N739_wire), .M1(M1[739:739]));

wire [7:0] ens0_layer0_N740_wire = {M0[13], M0[217], M0[354], M0[427], M0[504], M0[540], M0[578], M0[746]};
ens0_layer0_N740 ens0_layer0_N740_inst (.M0(ens0_layer0_N740_wire), .M1(M1[740:740]));

wire [7:0] ens0_layer0_N741_wire = {M0[51], M0[84], M0[123], M0[185], M0[409], M0[412], M0[492], M0[577]};
ens0_layer0_N741 ens0_layer0_N741_inst (.M0(ens0_layer0_N741_wire), .M1(M1[741:741]));

wire [7:0] ens0_layer0_N742_wire = {M0[11], M0[62], M0[90], M0[114], M0[149], M0[339], M0[354], M0[385]};
ens0_layer0_N742 ens0_layer0_N742_inst (.M0(ens0_layer0_N742_wire), .M1(M1[742:742]));

wire [7:0] ens0_layer0_N743_wire = {M0[54], M0[165], M0[237], M0[388], M0[416], M0[425], M0[567], M0[716]};
ens0_layer0_N743 ens0_layer0_N743_inst (.M0(ens0_layer0_N743_wire), .M1(M1[743:743]));

wire [7:0] ens0_layer0_N744_wire = {M0[87], M0[286], M0[326], M0[332], M0[530], M0[571], M0[608], M0[777]};
ens0_layer0_N744 ens0_layer0_N744_inst (.M0(ens0_layer0_N744_wire), .M1(M1[744:744]));

wire [7:0] ens0_layer0_N745_wire = {M0[21], M0[37], M0[116], M0[316], M0[325], M0[361], M0[596], M0[750]};
ens0_layer0_N745 ens0_layer0_N745_inst (.M0(ens0_layer0_N745_wire), .M1(M1[745:745]));

wire [7:0] ens0_layer0_N746_wire = {M0[94], M0[115], M0[223], M0[386], M0[391], M0[638], M0[658], M0[661]};
ens0_layer0_N746 ens0_layer0_N746_inst (.M0(ens0_layer0_N746_wire), .M1(M1[746:746]));

wire [7:0] ens0_layer0_N747_wire = {M0[13], M0[69], M0[171], M0[300], M0[472], M0[489], M0[693], M0[759]};
ens0_layer0_N747 ens0_layer0_N747_inst (.M0(ens0_layer0_N747_wire), .M1(M1[747:747]));

wire [7:0] ens0_layer0_N748_wire = {M0[191], M0[217], M0[250], M0[293], M0[426], M0[543], M0[654], M0[669]};
ens0_layer0_N748 ens0_layer0_N748_inst (.M0(ens0_layer0_N748_wire), .M1(M1[748:748]));

wire [7:0] ens0_layer0_N749_wire = {M0[51], M0[150], M0[180], M0[311], M0[468], M0[508], M0[693], M0[764]};
ens0_layer0_N749 ens0_layer0_N749_inst (.M0(ens0_layer0_N749_wire), .M1(M1[749:749]));

wire [7:0] ens0_layer0_N750_wire = {M0[57], M0[432], M0[441], M0[488], M0[599], M0[665], M0[742], M0[767]};
ens0_layer0_N750 ens0_layer0_N750_inst (.M0(ens0_layer0_N750_wire), .M1(M1[750:750]));

wire [7:0] ens0_layer0_N751_wire = {M0[207], M0[208], M0[251], M0[487], M0[488], M0[613], M0[663], M0[756]};
ens0_layer0_N751 ens0_layer0_N751_inst (.M0(ens0_layer0_N751_wire), .M1(M1[751:751]));

wire [7:0] ens0_layer0_N752_wire = {M0[222], M0[237], M0[318], M0[591], M0[621], M0[639], M0[764], M0[779]};
ens0_layer0_N752 ens0_layer0_N752_inst (.M0(ens0_layer0_N752_wire), .M1(M1[752:752]));

wire [7:0] ens0_layer0_N753_wire = {M0[102], M0[263], M0[315], M0[446], M0[529], M0[560], M0[567], M0[605]};
ens0_layer0_N753 ens0_layer0_N753_inst (.M0(ens0_layer0_N753_wire), .M1(M1[753:753]));

wire [7:0] ens0_layer0_N754_wire = {M0[82], M0[91], M0[122], M0[238], M0[375], M0[611], M0[619], M0[742]};
ens0_layer0_N754 ens0_layer0_N754_inst (.M0(ens0_layer0_N754_wire), .M1(M1[754:754]));

wire [7:0] ens0_layer0_N755_wire = {M0[133], M0[142], M0[195], M0[211], M0[230], M0[378], M0[545], M0[672]};
ens0_layer0_N755 ens0_layer0_N755_inst (.M0(ens0_layer0_N755_wire), .M1(M1[755:755]));

wire [7:0] ens0_layer0_N756_wire = {M0[9], M0[164], M0[219], M0[354], M0[408], M0[557], M0[564], M0[700]};
ens0_layer0_N756 ens0_layer0_N756_inst (.M0(ens0_layer0_N756_wire), .M1(M1[756:756]));

wire [7:0] ens0_layer0_N757_wire = {M0[141], M0[148], M0[215], M0[256], M0[565], M0[603], M0[608], M0[636]};
ens0_layer0_N757 ens0_layer0_N757_inst (.M0(ens0_layer0_N757_wire), .M1(M1[757:757]));

wire [7:0] ens0_layer0_N758_wire = {M0[0], M0[97], M0[114], M0[137], M0[199], M0[591], M0[634], M0[664]};
ens0_layer0_N758 ens0_layer0_N758_inst (.M0(ens0_layer0_N758_wire), .M1(M1[758:758]));

wire [7:0] ens0_layer0_N759_wire = {M0[34], M0[111], M0[200], M0[367], M0[514], M0[553], M0[657], M0[762]};
ens0_layer0_N759 ens0_layer0_N759_inst (.M0(ens0_layer0_N759_wire), .M1(M1[759:759]));

wire [7:0] ens0_layer0_N760_wire = {M0[99], M0[106], M0[140], M0[300], M0[316], M0[322], M0[398], M0[648]};
ens0_layer0_N760 ens0_layer0_N760_inst (.M0(ens0_layer0_N760_wire), .M1(M1[760:760]));

wire [7:0] ens0_layer0_N761_wire = {M0[140], M0[169], M0[179], M0[241], M0[417], M0[466], M0[653], M0[773]};
ens0_layer0_N761 ens0_layer0_N761_inst (.M0(ens0_layer0_N761_wire), .M1(M1[761:761]));

wire [7:0] ens0_layer0_N762_wire = {M0[18], M0[29], M0[66], M0[347], M0[372], M0[485], M0[565], M0[627]};
ens0_layer0_N762 ens0_layer0_N762_inst (.M0(ens0_layer0_N762_wire), .M1(M1[762:762]));

wire [7:0] ens0_layer0_N763_wire = {M0[224], M0[302], M0[372], M0[377], M0[437], M0[627], M0[760], M0[779]};
ens0_layer0_N763 ens0_layer0_N763_inst (.M0(ens0_layer0_N763_wire), .M1(M1[763:763]));

wire [7:0] ens0_layer0_N764_wire = {M0[12], M0[106], M0[245], M0[520], M0[549], M0[577], M0[718], M0[741]};
ens0_layer0_N764 ens0_layer0_N764_inst (.M0(ens0_layer0_N764_wire), .M1(M1[764:764]));

wire [7:0] ens0_layer0_N765_wire = {M0[162], M0[197], M0[205], M0[308], M0[328], M0[364], M0[391], M0[509]};
ens0_layer0_N765 ens0_layer0_N765_inst (.M0(ens0_layer0_N765_wire), .M1(M1[765:765]));

wire [7:0] ens0_layer0_N766_wire = {M0[122], M0[250], M0[285], M0[440], M0[626], M0[727], M0[756], M0[775]};
ens0_layer0_N766 ens0_layer0_N766_inst (.M0(ens0_layer0_N766_wire), .M1(M1[766:766]));

wire [7:0] ens0_layer0_N767_wire = {M0[123], M0[138], M0[318], M0[463], M0[502], M0[642], M0[671], M0[718]};
ens0_layer0_N767 ens0_layer0_N767_inst (.M0(ens0_layer0_N767_wire), .M1(M1[767:767]));

wire [7:0] ens0_layer0_N768_wire = {M0[25], M0[34], M0[289], M0[373], M0[445], M0[570], M0[589], M0[718]};
ens0_layer0_N768 ens0_layer0_N768_inst (.M0(ens0_layer0_N768_wire), .M1(M1[768:768]));

wire [7:0] ens0_layer0_N769_wire = {M0[92], M0[136], M0[159], M0[202], M0[447], M0[449], M0[458], M0[704]};
ens0_layer0_N769 ens0_layer0_N769_inst (.M0(ens0_layer0_N769_wire), .M1(M1[769:769]));

wire [7:0] ens0_layer0_N770_wire = {M0[22], M0[229], M0[296], M0[345], M0[431], M0[465], M0[547], M0[700]};
ens0_layer0_N770 ens0_layer0_N770_inst (.M0(ens0_layer0_N770_wire), .M1(M1[770:770]));

wire [7:0] ens0_layer0_N771_wire = {M0[212], M0[224], M0[240], M0[324], M0[447], M0[611], M0[715], M0[751]};
ens0_layer0_N771 ens0_layer0_N771_inst (.M0(ens0_layer0_N771_wire), .M1(M1[771:771]));

wire [7:0] ens0_layer0_N772_wire = {M0[67], M0[249], M0[276], M0[354], M0[467], M0[608], M0[649], M0[650]};
ens0_layer0_N772 ens0_layer0_N772_inst (.M0(ens0_layer0_N772_wire), .M1(M1[772:772]));

wire [7:0] ens0_layer0_N773_wire = {M0[7], M0[225], M0[394], M0[484], M0[493], M0[515], M0[644], M0[690]};
ens0_layer0_N773 ens0_layer0_N773_inst (.M0(ens0_layer0_N773_wire), .M1(M1[773:773]));

wire [7:0] ens0_layer0_N774_wire = {M0[130], M0[145], M0[301], M0[370], M0[425], M0[541], M0[583], M0[658]};
ens0_layer0_N774 ens0_layer0_N774_inst (.M0(ens0_layer0_N774_wire), .M1(M1[774:774]));

wire [7:0] ens0_layer0_N775_wire = {M0[39], M0[48], M0[90], M0[93], M0[99], M0[342], M0[384], M0[731]};
ens0_layer0_N775 ens0_layer0_N775_inst (.M0(ens0_layer0_N775_wire), .M1(M1[775:775]));

wire [7:0] ens0_layer0_N776_wire = {M0[29], M0[280], M0[329], M0[423], M0[476], M0[539], M0[605], M0[683]};
ens0_layer0_N776 ens0_layer0_N776_inst (.M0(ens0_layer0_N776_wire), .M1(M1[776:776]));

wire [7:0] ens0_layer0_N777_wire = {M0[107], M0[160], M0[172], M0[454], M0[494], M0[504], M0[612], M0[757]};
ens0_layer0_N777 ens0_layer0_N777_inst (.M0(ens0_layer0_N777_wire), .M1(M1[777:777]));

wire [7:0] ens0_layer0_N778_wire = {M0[29], M0[82], M0[417], M0[502], M0[607], M0[759], M0[771], M0[773]};
ens0_layer0_N778 ens0_layer0_N778_inst (.M0(ens0_layer0_N778_wire), .M1(M1[778:778]));

wire [7:0] ens0_layer0_N779_wire = {M0[197], M0[325], M0[396], M0[486], M0[495], M0[618], M0[634], M0[755]};
ens0_layer0_N779 ens0_layer0_N779_inst (.M0(ens0_layer0_N779_wire), .M1(M1[779:779]));

wire [7:0] ens0_layer0_N780_wire = {M0[104], M0[115], M0[139], M0[206], M0[265], M0[350], M0[533], M0[746]};
ens0_layer0_N780 ens0_layer0_N780_inst (.M0(ens0_layer0_N780_wire), .M1(M1[780:780]));

wire [7:0] ens0_layer0_N781_wire = {M0[37], M0[266], M0[289], M0[533], M0[593], M0[619], M0[655], M0[741]};
ens0_layer0_N781 ens0_layer0_N781_inst (.M0(ens0_layer0_N781_wire), .M1(M1[781:781]));

wire [7:0] ens0_layer0_N782_wire = {M0[22], M0[92], M0[145], M0[188], M0[217], M0[526], M0[701], M0[775]};
ens0_layer0_N782 ens0_layer0_N782_inst (.M0(ens0_layer0_N782_wire), .M1(M1[782:782]));

wire [7:0] ens0_layer0_N783_wire = {M0[46], M0[79], M0[300], M0[362], M0[567], M0[585], M0[630], M0[715]};
ens0_layer0_N783 ens0_layer0_N783_inst (.M0(ens0_layer0_N783_wire), .M1(M1[783:783]));

wire [7:0] ens0_layer0_N784_wire = {M0[16], M0[87], M0[122], M0[171], M0[234], M0[247], M0[333], M0[742]};
ens0_layer0_N784 ens0_layer0_N784_inst (.M0(ens0_layer0_N784_wire), .M1(M1[784:784]));

wire [7:0] ens0_layer0_N785_wire = {M0[81], M0[87], M0[115], M0[205], M0[368], M0[605], M0[611], M0[669]};
ens0_layer0_N785 ens0_layer0_N785_inst (.M0(ens0_layer0_N785_wire), .M1(M1[785:785]));

wire [7:0] ens0_layer0_N786_wire = {M0[143], M0[181], M0[224], M0[356], M0[407], M0[450], M0[547], M0[687]};
ens0_layer0_N786 ens0_layer0_N786_inst (.M0(ens0_layer0_N786_wire), .M1(M1[786:786]));

wire [7:0] ens0_layer0_N787_wire = {M0[124], M0[246], M0[254], M0[418], M0[439], M0[454], M0[665], M0[730]};
ens0_layer0_N787 ens0_layer0_N787_inst (.M0(ens0_layer0_N787_wire), .M1(M1[787:787]));

wire [7:0] ens0_layer0_N788_wire = {M0[15], M0[118], M0[188], M0[222], M0[376], M0[410], M0[511], M0[570]};
ens0_layer0_N788 ens0_layer0_N788_inst (.M0(ens0_layer0_N788_wire), .M1(M1[788:788]));

wire [7:0] ens0_layer0_N789_wire = {M0[81], M0[224], M0[289], M0[407], M0[486], M0[521], M0[735], M0[772]};
ens0_layer0_N789 ens0_layer0_N789_inst (.M0(ens0_layer0_N789_wire), .M1(M1[789:789]));

wire [7:0] ens0_layer0_N790_wire = {M0[54], M0[118], M0[253], M0[296], M0[329], M0[406], M0[461], M0[507]};
ens0_layer0_N790 ens0_layer0_N790_inst (.M0(ens0_layer0_N790_wire), .M1(M1[790:790]));

wire [7:0] ens0_layer0_N791_wire = {M0[213], M0[280], M0[443], M0[450], M0[564], M0[609], M0[666], M0[772]};
ens0_layer0_N791 ens0_layer0_N791_inst (.M0(ens0_layer0_N791_wire), .M1(M1[791:791]));

wire [7:0] ens0_layer0_N792_wire = {M0[264], M0[329], M0[404], M0[503], M0[529], M0[650], M0[714], M0[768]};
ens0_layer0_N792 ens0_layer0_N792_inst (.M0(ens0_layer0_N792_wire), .M1(M1[792:792]));

wire [7:0] ens0_layer0_N793_wire = {M0[48], M0[423], M0[495], M0[615], M0[622], M0[688], M0[752], M0[778]};
ens0_layer0_N793 ens0_layer0_N793_inst (.M0(ens0_layer0_N793_wire), .M1(M1[793:793]));

wire [7:0] ens0_layer0_N794_wire = {M0[151], M0[219], M0[437], M0[453], M0[557], M0[665], M0[737], M0[783]};
ens0_layer0_N794 ens0_layer0_N794_inst (.M0(ens0_layer0_N794_wire), .M1(M1[794:794]));

wire [7:0] ens0_layer0_N795_wire = {M0[109], M0[110], M0[203], M0[423], M0[510], M0[563], M0[609], M0[733]};
ens0_layer0_N795 ens0_layer0_N795_inst (.M0(ens0_layer0_N795_wire), .M1(M1[795:795]));

wire [7:0] ens0_layer0_N796_wire = {M0[85], M0[443], M0[489], M0[574], M0[594], M0[603], M0[721], M0[774]};
ens0_layer0_N796 ens0_layer0_N796_inst (.M0(ens0_layer0_N796_wire), .M1(M1[796:796]));

wire [7:0] ens0_layer0_N797_wire = {M0[20], M0[90], M0[218], M0[458], M0[577], M0[588], M0[700], M0[774]};
ens0_layer0_N797 ens0_layer0_N797_inst (.M0(ens0_layer0_N797_wire), .M1(M1[797:797]));

wire [7:0] ens0_layer0_N798_wire = {M0[84], M0[122], M0[263], M0[353], M0[412], M0[474], M0[638], M0[715]};
ens0_layer0_N798 ens0_layer0_N798_inst (.M0(ens0_layer0_N798_wire), .M1(M1[798:798]));

wire [7:0] ens0_layer0_N799_wire = {M0[106], M0[129], M0[369], M0[371], M0[404], M0[578], M0[683], M0[726]};
ens0_layer0_N799 ens0_layer0_N799_inst (.M0(ens0_layer0_N799_wire), .M1(M1[799:799]));

wire [7:0] ens0_layer0_N800_wire = {M0[20], M0[62], M0[167], M0[365], M0[512], M0[595], M0[665], M0[781]};
ens0_layer0_N800 ens0_layer0_N800_inst (.M0(ens0_layer0_N800_wire), .M1(M1[800:800]));

wire [7:0] ens0_layer0_N801_wire = {M0[46], M0[70], M0[89], M0[212], M0[295], M0[350], M0[369], M0[467]};
ens0_layer0_N801 ens0_layer0_N801_inst (.M0(ens0_layer0_N801_wire), .M1(M1[801:801]));

wire [7:0] ens0_layer0_N802_wire = {M0[75], M0[106], M0[140], M0[148], M0[264], M0[669], M0[747], M0[775]};
ens0_layer0_N802 ens0_layer0_N802_inst (.M0(ens0_layer0_N802_wire), .M1(M1[802:802]));

wire [7:0] ens0_layer0_N803_wire = {M0[3], M0[31], M0[69], M0[114], M0[141], M0[350], M0[435], M0[480]};
ens0_layer0_N803 ens0_layer0_N803_inst (.M0(ens0_layer0_N803_wire), .M1(M1[803:803]));

wire [7:0] ens0_layer0_N804_wire = {M0[64], M0[118], M0[124], M0[139], M0[150], M0[214], M0[326], M0[772]};
ens0_layer0_N804 ens0_layer0_N804_inst (.M0(ens0_layer0_N804_wire), .M1(M1[804:804]));

wire [7:0] ens0_layer0_N805_wire = {M0[47], M0[97], M0[178], M0[242], M0[334], M0[357], M0[692], M0[759]};
ens0_layer0_N805 ens0_layer0_N805_inst (.M0(ens0_layer0_N805_wire), .M1(M1[805:805]));

wire [7:0] ens0_layer0_N806_wire = {M0[64], M0[169], M0[336], M0[449], M0[557], M0[589], M0[718], M0[745]};
ens0_layer0_N806 ens0_layer0_N806_inst (.M0(ens0_layer0_N806_wire), .M1(M1[806:806]));

wire [7:0] ens0_layer0_N807_wire = {M0[30], M0[122], M0[253], M0[430], M0[468], M0[564], M0[689], M0[697]};
ens0_layer0_N807 ens0_layer0_N807_inst (.M0(ens0_layer0_N807_wire), .M1(M1[807:807]));

wire [7:0] ens0_layer0_N808_wire = {M0[74], M0[145], M0[212], M0[261], M0[369], M0[530], M0[579], M0[605]};
ens0_layer0_N808 ens0_layer0_N808_inst (.M0(ens0_layer0_N808_wire), .M1(M1[808:808]));

wire [7:0] ens0_layer0_N809_wire = {M0[24], M0[186], M0[316], M0[322], M0[332], M0[442], M0[453], M0[544]};
ens0_layer0_N809 ens0_layer0_N809_inst (.M0(ens0_layer0_N809_wire), .M1(M1[809:809]));

wire [7:0] ens0_layer0_N810_wire = {M0[139], M0[166], M0[175], M0[203], M0[499], M0[633], M0[707], M0[730]};
ens0_layer0_N810 ens0_layer0_N810_inst (.M0(ens0_layer0_N810_wire), .M1(M1[810:810]));

wire [7:0] ens0_layer0_N811_wire = {M0[103], M0[144], M0[290], M0[347], M0[443], M0[527], M0[704], M0[759]};
ens0_layer0_N811 ens0_layer0_N811_inst (.M0(ens0_layer0_N811_wire), .M1(M1[811:811]));

wire [7:0] ens0_layer0_N812_wire = {M0[40], M0[70], M0[123], M0[124], M0[157], M0[507], M0[539], M0[647]};
ens0_layer0_N812 ens0_layer0_N812_inst (.M0(ens0_layer0_N812_wire), .M1(M1[812:812]));

wire [7:0] ens0_layer0_N813_wire = {M0[22], M0[95], M0[306], M0[333], M0[335], M0[405], M0[498], M0[750]};
ens0_layer0_N813 ens0_layer0_N813_inst (.M0(ens0_layer0_N813_wire), .M1(M1[813:813]));

wire [7:0] ens0_layer0_N814_wire = {M0[20], M0[45], M0[155], M0[378], M0[479], M0[490], M0[511], M0[596]};
ens0_layer0_N814 ens0_layer0_N814_inst (.M0(ens0_layer0_N814_wire), .M1(M1[814:814]));

wire [7:0] ens0_layer0_N815_wire = {M0[269], M0[281], M0[334], M0[387], M0[497], M0[507], M0[688], M0[728]};
ens0_layer0_N815 ens0_layer0_N815_inst (.M0(ens0_layer0_N815_wire), .M1(M1[815:815]));

wire [7:0] ens0_layer0_N816_wire = {M0[248], M0[256], M0[264], M0[333], M0[506], M0[515], M0[552], M0[700]};
ens0_layer0_N816 ens0_layer0_N816_inst (.M0(ens0_layer0_N816_wire), .M1(M1[816:816]));

wire [7:0] ens0_layer0_N817_wire = {M0[0], M0[96], M0[245], M0[350], M0[408], M0[476], M0[529], M0[584]};
ens0_layer0_N817 ens0_layer0_N817_inst (.M0(ens0_layer0_N817_wire), .M1(M1[817:817]));

wire [7:0] ens0_layer0_N818_wire = {M0[72], M0[191], M0[231], M0[338], M0[391], M0[471], M0[588], M0[603]};
ens0_layer0_N818 ens0_layer0_N818_inst (.M0(ens0_layer0_N818_wire), .M1(M1[818:818]));

wire [7:0] ens0_layer0_N819_wire = {M0[70], M0[95], M0[191], M0[198], M0[538], M0[576], M0[772], M0[780]};
ens0_layer0_N819 ens0_layer0_N819_inst (.M0(ens0_layer0_N819_wire), .M1(M1[819:819]));

wire [7:0] ens0_layer0_N820_wire = {M0[47], M0[48], M0[81], M0[118], M0[226], M0[283], M0[592], M0[733]};
ens0_layer0_N820 ens0_layer0_N820_inst (.M0(ens0_layer0_N820_wire), .M1(M1[820:820]));

wire [7:0] ens0_layer0_N821_wire = {M0[144], M0[255], M0[308], M0[343], M0[414], M0[571], M0[719], M0[745]};
ens0_layer0_N821 ens0_layer0_N821_inst (.M0(ens0_layer0_N821_wire), .M1(M1[821:821]));

wire [7:0] ens0_layer0_N822_wire = {M0[18], M0[32], M0[92], M0[102], M0[175], M0[454], M0[466], M0[516]};
ens0_layer0_N822 ens0_layer0_N822_inst (.M0(ens0_layer0_N822_wire), .M1(M1[822:822]));

wire [7:0] ens0_layer0_N823_wire = {M0[129], M0[170], M0[211], M0[302], M0[305], M0[381], M0[620], M0[741]};
ens0_layer0_N823 ens0_layer0_N823_inst (.M0(ens0_layer0_N823_wire), .M1(M1[823:823]));

wire [7:0] ens0_layer0_N824_wire = {M0[15], M0[36], M0[115], M0[151], M0[215], M0[569], M0[633], M0[650]};
ens0_layer0_N824 ens0_layer0_N824_inst (.M0(ens0_layer0_N824_wire), .M1(M1[824:824]));

wire [7:0] ens0_layer0_N825_wire = {M0[144], M0[176], M0[231], M0[457], M0[560], M0[639], M0[705], M0[739]};
ens0_layer0_N825 ens0_layer0_N825_inst (.M0(ens0_layer0_N825_wire), .M1(M1[825:825]));

wire [7:0] ens0_layer0_N826_wire = {M0[13], M0[55], M0[58], M0[168], M0[390], M0[451], M0[474], M0[682]};
ens0_layer0_N826 ens0_layer0_N826_inst (.M0(ens0_layer0_N826_wire), .M1(M1[826:826]));

wire [7:0] ens0_layer0_N827_wire = {M0[55], M0[155], M0[201], M0[243], M0[349], M0[352], M0[535], M0[575]};
ens0_layer0_N827 ens0_layer0_N827_inst (.M0(ens0_layer0_N827_wire), .M1(M1[827:827]));

wire [7:0] ens0_layer0_N828_wire = {M0[208], M0[446], M0[465], M0[470], M0[544], M0[611], M0[664], M0[783]};
ens0_layer0_N828 ens0_layer0_N828_inst (.M0(ens0_layer0_N828_wire), .M1(M1[828:828]));

wire [7:0] ens0_layer0_N829_wire = {M0[23], M0[58], M0[342], M0[424], M0[425], M0[471], M0[539], M0[595]};
ens0_layer0_N829 ens0_layer0_N829_inst (.M0(ens0_layer0_N829_wire), .M1(M1[829:829]));

wire [7:0] ens0_layer0_N830_wire = {M0[85], M0[156], M0[388], M0[420], M0[474], M0[616], M0[631], M0[737]};
ens0_layer0_N830 ens0_layer0_N830_inst (.M0(ens0_layer0_N830_wire), .M1(M1[830:830]));

wire [7:0] ens0_layer0_N831_wire = {M0[21], M0[303], M0[351], M0[505], M0[537], M0[569], M0[607], M0[713]};
ens0_layer0_N831 ens0_layer0_N831_inst (.M0(ens0_layer0_N831_wire), .M1(M1[831:831]));

wire [7:0] ens0_layer0_N832_wire = {M0[60], M0[103], M0[148], M0[149], M0[173], M0[272], M0[602], M0[719]};
ens0_layer0_N832 ens0_layer0_N832_inst (.M0(ens0_layer0_N832_wire), .M1(M1[832:832]));

wire [7:0] ens0_layer0_N833_wire = {M0[31], M0[301], M0[328], M0[355], M0[514], M0[528], M0[536], M0[712]};
ens0_layer0_N833 ens0_layer0_N833_inst (.M0(ens0_layer0_N833_wire), .M1(M1[833:833]));

wire [7:0] ens0_layer0_N834_wire = {M0[104], M0[150], M0[152], M0[539], M0[619], M0[624], M0[704], M0[710]};
ens0_layer0_N834 ens0_layer0_N834_inst (.M0(ens0_layer0_N834_wire), .M1(M1[834:834]));

wire [7:0] ens0_layer0_N835_wire = {M0[57], M0[65], M0[81], M0[371], M0[428], M0[468], M0[498], M0[551]};
ens0_layer0_N835 ens0_layer0_N835_inst (.M0(ens0_layer0_N835_wire), .M1(M1[835:835]));

wire [7:0] ens0_layer0_N836_wire = {M0[8], M0[132], M0[261], M0[583], M0[736], M0[737], M0[743], M0[745]};
ens0_layer0_N836 ens0_layer0_N836_inst (.M0(ens0_layer0_N836_wire), .M1(M1[836:836]));

wire [7:0] ens0_layer0_N837_wire = {M0[14], M0[99], M0[175], M0[483], M0[507], M0[579], M0[690], M0[762]};
ens0_layer0_N837 ens0_layer0_N837_inst (.M0(ens0_layer0_N837_wire), .M1(M1[837:837]));

wire [7:0] ens0_layer0_N838_wire = {M0[146], M0[234], M0[266], M0[385], M0[634], M0[648], M0[695], M0[718]};
ens0_layer0_N838 ens0_layer0_N838_inst (.M0(ens0_layer0_N838_wire), .M1(M1[838:838]));

wire [7:0] ens0_layer0_N839_wire = {M0[5], M0[101], M0[151], M0[188], M0[409], M0[442], M0[671], M0[732]};
ens0_layer0_N839 ens0_layer0_N839_inst (.M0(ens0_layer0_N839_wire), .M1(M1[839:839]));

wire [7:0] ens0_layer0_N840_wire = {M0[121], M0[151], M0[188], M0[250], M0[392], M0[478], M0[695], M0[732]};
ens0_layer0_N840 ens0_layer0_N840_inst (.M0(ens0_layer0_N840_wire), .M1(M1[840:840]));

wire [7:0] ens0_layer0_N841_wire = {M0[161], M0[215], M0[221], M0[229], M0[240], M0[318], M0[369], M0[601]};
ens0_layer0_N841 ens0_layer0_N841_inst (.M0(ens0_layer0_N841_wire), .M1(M1[841:841]));

wire [7:0] ens0_layer0_N842_wire = {M0[112], M0[234], M0[304], M0[405], M0[448], M0[534], M0[564], M0[772]};
ens0_layer0_N842 ens0_layer0_N842_inst (.M0(ens0_layer0_N842_wire), .M1(M1[842:842]));

wire [7:0] ens0_layer0_N843_wire = {M0[34], M0[251], M0[298], M0[357], M0[441], M0[458], M0[486], M0[751]};
ens0_layer0_N843 ens0_layer0_N843_inst (.M0(ens0_layer0_N843_wire), .M1(M1[843:843]));

wire [7:0] ens0_layer0_N844_wire = {M0[123], M0[317], M0[374], M0[475], M0[558], M0[690], M0[747], M0[763]};
ens0_layer0_N844 ens0_layer0_N844_inst (.M0(ens0_layer0_N844_wire), .M1(M1[844:844]));

wire [7:0] ens0_layer0_N845_wire = {M0[41], M0[66], M0[125], M0[242], M0[345], M0[360], M0[437], M0[690]};
ens0_layer0_N845 ens0_layer0_N845_inst (.M0(ens0_layer0_N845_wire), .M1(M1[845:845]));

wire [7:0] ens0_layer0_N846_wire = {M0[235], M0[261], M0[269], M0[291], M0[334], M0[647], M0[648], M0[700]};
ens0_layer0_N846 ens0_layer0_N846_inst (.M0(ens0_layer0_N846_wire), .M1(M1[846:846]));

wire [7:0] ens0_layer0_N847_wire = {M0[148], M0[162], M0[201], M0[218], M0[543], M0[696], M0[703], M0[750]};
ens0_layer0_N847 ens0_layer0_N847_inst (.M0(ens0_layer0_N847_wire), .M1(M1[847:847]));

wire [7:0] ens0_layer0_N848_wire = {M0[90], M0[243], M0[355], M0[365], M0[527], M0[533], M0[583], M0[710]};
ens0_layer0_N848 ens0_layer0_N848_inst (.M0(ens0_layer0_N848_wire), .M1(M1[848:848]));

wire [7:0] ens0_layer0_N849_wire = {M0[152], M0[203], M0[370], M0[464], M0[614], M0[641], M0[693], M0[781]};
ens0_layer0_N849 ens0_layer0_N849_inst (.M0(ens0_layer0_N849_wire), .M1(M1[849:849]));

wire [7:0] ens0_layer0_N850_wire = {M0[64], M0[121], M0[327], M0[359], M0[372], M0[419], M0[651], M0[664]};
ens0_layer0_N850 ens0_layer0_N850_inst (.M0(ens0_layer0_N850_wire), .M1(M1[850:850]));

wire [7:0] ens0_layer0_N851_wire = {M0[211], M0[248], M0[345], M0[378], M0[493], M0[528], M0[555], M0[764]};
ens0_layer0_N851 ens0_layer0_N851_inst (.M0(ens0_layer0_N851_wire), .M1(M1[851:851]));

wire [7:0] ens0_layer0_N852_wire = {M0[29], M0[108], M0[171], M0[237], M0[269], M0[411], M0[510], M0[597]};
ens0_layer0_N852 ens0_layer0_N852_inst (.M0(ens0_layer0_N852_wire), .M1(M1[852:852]));

wire [7:0] ens0_layer0_N853_wire = {M0[75], M0[77], M0[298], M0[525], M0[614], M0[664], M0[722], M0[735]};
ens0_layer0_N853 ens0_layer0_N853_inst (.M0(ens0_layer0_N853_wire), .M1(M1[853:853]));

wire [7:0] ens0_layer0_N854_wire = {M0[11], M0[120], M0[134], M0[217], M0[295], M0[486], M0[642], M0[737]};
ens0_layer0_N854 ens0_layer0_N854_inst (.M0(ens0_layer0_N854_wire), .M1(M1[854:854]));

wire [7:0] ens0_layer0_N855_wire = {M0[124], M0[153], M0[317], M0[392], M0[465], M0[520], M0[532], M0[656]};
ens0_layer0_N855 ens0_layer0_N855_inst (.M0(ens0_layer0_N855_wire), .M1(M1[855:855]));

wire [7:0] ens0_layer0_N856_wire = {M0[160], M0[429], M0[452], M0[489], M0[553], M0[556], M0[569], M0[667]};
ens0_layer0_N856 ens0_layer0_N856_inst (.M0(ens0_layer0_N856_wire), .M1(M1[856:856]));

wire [7:0] ens0_layer0_N857_wire = {M0[33], M0[72], M0[112], M0[373], M0[429], M0[439], M0[535], M0[742]};
ens0_layer0_N857 ens0_layer0_N857_inst (.M0(ens0_layer0_N857_wire), .M1(M1[857:857]));

wire [7:0] ens0_layer0_N858_wire = {M0[509], M0[550], M0[558], M0[585], M0[617], M0[694], M0[717], M0[728]};
ens0_layer0_N858 ens0_layer0_N858_inst (.M0(ens0_layer0_N858_wire), .M1(M1[858:858]));

wire [7:0] ens0_layer0_N859_wire = {M0[268], M0[432], M0[448], M0[501], M0[516], M0[629], M0[647], M0[753]};
ens0_layer0_N859 ens0_layer0_N859_inst (.M0(ens0_layer0_N859_wire), .M1(M1[859:859]));

wire [7:0] ens0_layer0_N860_wire = {M0[17], M0[204], M0[236], M0[252], M0[340], M0[354], M0[597], M0[741]};
ens0_layer0_N860 ens0_layer0_N860_inst (.M0(ens0_layer0_N860_wire), .M1(M1[860:860]));

wire [7:0] ens0_layer0_N861_wire = {M0[102], M0[389], M0[461], M0[540], M0[545], M0[638], M0[671], M0[695]};
ens0_layer0_N861 ens0_layer0_N861_inst (.M0(ens0_layer0_N861_wire), .M1(M1[861:861]));

wire [7:0] ens0_layer0_N862_wire = {M0[10], M0[134], M0[225], M0[250], M0[504], M0[632], M0[701], M0[744]};
ens0_layer0_N862 ens0_layer0_N862_inst (.M0(ens0_layer0_N862_wire), .M1(M1[862:862]));

wire [7:0] ens0_layer0_N863_wire = {M0[94], M0[170], M0[372], M0[373], M0[439], M0[581], M0[694], M0[715]};
ens0_layer0_N863 ens0_layer0_N863_inst (.M0(ens0_layer0_N863_wire), .M1(M1[863:863]));

wire [7:0] ens0_layer0_N864_wire = {M0[8], M0[270], M0[344], M0[445], M0[535], M0[601], M0[714], M0[753]};
ens0_layer0_N864 ens0_layer0_N864_inst (.M0(ens0_layer0_N864_wire), .M1(M1[864:864]));

wire [7:0] ens0_layer0_N865_wire = {M0[1], M0[101], M0[123], M0[125], M0[370], M0[616], M0[625], M0[753]};
ens0_layer0_N865 ens0_layer0_N865_inst (.M0(ens0_layer0_N865_wire), .M1(M1[865:865]));

wire [7:0] ens0_layer0_N866_wire = {M0[84], M0[153], M0[193], M0[415], M0[500], M0[607], M0[692], M0[768]};
ens0_layer0_N866 ens0_layer0_N866_inst (.M0(ens0_layer0_N866_wire), .M1(M1[866:866]));

wire [7:0] ens0_layer0_N867_wire = {M0[16], M0[230], M0[383], M0[414], M0[437], M0[564], M0[585], M0[705]};
ens0_layer0_N867 ens0_layer0_N867_inst (.M0(ens0_layer0_N867_wire), .M1(M1[867:867]));

wire [7:0] ens0_layer0_N868_wire = {M0[17], M0[204], M0[345], M0[479], M0[590], M0[629], M0[697], M0[698]};
ens0_layer0_N868 ens0_layer0_N868_inst (.M0(ens0_layer0_N868_wire), .M1(M1[868:868]));

wire [7:0] ens0_layer0_N869_wire = {M0[146], M0[236], M0[286], M0[327], M0[377], M0[400], M0[444], M0[547]};
ens0_layer0_N869 ens0_layer0_N869_inst (.M0(ens0_layer0_N869_wire), .M1(M1[869:869]));

wire [7:0] ens0_layer0_N870_wire = {M0[99], M0[173], M0[208], M0[377], M0[669], M0[735], M0[738], M0[749]};
ens0_layer0_N870 ens0_layer0_N870_inst (.M0(ens0_layer0_N870_wire), .M1(M1[870:870]));

wire [7:0] ens0_layer0_N871_wire = {M0[127], M0[207], M0[273], M0[292], M0[455], M0[618], M0[665], M0[683]};
ens0_layer0_N871 ens0_layer0_N871_inst (.M0(ens0_layer0_N871_wire), .M1(M1[871:871]));

wire [7:0] ens0_layer0_N872_wire = {M0[12], M0[123], M0[341], M0[365], M0[449], M0[535], M0[762], M0[780]};
ens0_layer0_N872 ens0_layer0_N872_inst (.M0(ens0_layer0_N872_wire), .M1(M1[872:872]));

wire [7:0] ens0_layer0_N873_wire = {M0[95], M0[176], M0[493], M0[513], M0[580], M0[635], M0[648], M0[751]};
ens0_layer0_N873 ens0_layer0_N873_inst (.M0(ens0_layer0_N873_wire), .M1(M1[873:873]));

wire [7:0] ens0_layer0_N874_wire = {M0[18], M0[90], M0[160], M0[168], M0[292], M0[431], M0[438], M0[738]};
ens0_layer0_N874 ens0_layer0_N874_inst (.M0(ens0_layer0_N874_wire), .M1(M1[874:874]));

wire [7:0] ens0_layer0_N875_wire = {M0[42], M0[176], M0[452], M0[543], M0[606], M0[646], M0[722], M0[734]};
ens0_layer0_N875 ens0_layer0_N875_inst (.M0(ens0_layer0_N875_wire), .M1(M1[875:875]));

wire [7:0] ens0_layer0_N876_wire = {M0[77], M0[79], M0[172], M0[195], M0[211], M0[301], M0[369], M0[493]};
ens0_layer0_N876 ens0_layer0_N876_inst (.M0(ens0_layer0_N876_wire), .M1(M1[876:876]));

wire [7:0] ens0_layer0_N877_wire = {M0[137], M0[350], M0[355], M0[456], M0[473], M0[517], M0[711], M0[727]};
ens0_layer0_N877 ens0_layer0_N877_inst (.M0(ens0_layer0_N877_wire), .M1(M1[877:877]));

wire [7:0] ens0_layer0_N878_wire = {M0[24], M0[59], M0[66], M0[126], M0[189], M0[468], M0[522], M0[767]};
ens0_layer0_N878 ens0_layer0_N878_inst (.M0(ens0_layer0_N878_wire), .M1(M1[878:878]));

wire [7:0] ens0_layer0_N879_wire = {M0[191], M0[242], M0[404], M0[431], M0[598], M0[623], M0[713], M0[759]};
ens0_layer0_N879 ens0_layer0_N879_inst (.M0(ens0_layer0_N879_wire), .M1(M1[879:879]));

wire [7:0] ens0_layer0_N880_wire = {M0[37], M0[46], M0[60], M0[76], M0[103], M0[148], M0[310], M0[419]};
ens0_layer0_N880 ens0_layer0_N880_inst (.M0(ens0_layer0_N880_wire), .M1(M1[880:880]));

wire [7:0] ens0_layer0_N881_wire = {M0[58], M0[354], M0[401], M0[472], M0[608], M0[734], M0[756], M0[762]};
ens0_layer0_N881 ens0_layer0_N881_inst (.M0(ens0_layer0_N881_wire), .M1(M1[881:881]));

wire [7:0] ens0_layer0_N882_wire = {M0[82], M0[152], M0[156], M0[159], M0[181], M0[363], M0[404], M0[500]};
ens0_layer0_N882 ens0_layer0_N882_inst (.M0(ens0_layer0_N882_wire), .M1(M1[882:882]));

wire [7:0] ens0_layer0_N883_wire = {M0[114], M0[278], M0[285], M0[318], M0[366], M0[434], M0[605], M0[724]};
ens0_layer0_N883 ens0_layer0_N883_inst (.M0(ens0_layer0_N883_wire), .M1(M1[883:883]));

wire [7:0] ens0_layer0_N884_wire = {M0[45], M0[158], M0[221], M0[419], M0[528], M0[579], M0[587], M0[684]};
ens0_layer0_N884 ens0_layer0_N884_inst (.M0(ens0_layer0_N884_wire), .M1(M1[884:884]));

wire [7:0] ens0_layer0_N885_wire = {M0[9], M0[37], M0[75], M0[228], M0[346], M0[507], M0[531], M0[671]};
ens0_layer0_N885 ens0_layer0_N885_inst (.M0(ens0_layer0_N885_wire), .M1(M1[885:885]));

wire [7:0] ens0_layer0_N886_wire = {M0[145], M0[230], M0[507], M0[570], M0[670], M0[684], M0[725], M0[773]};
ens0_layer0_N886 ens0_layer0_N886_inst (.M0(ens0_layer0_N886_wire), .M1(M1[886:886]));

wire [7:0] ens0_layer0_N887_wire = {M0[9], M0[86], M0[249], M0[489], M0[516], M0[556], M0[622], M0[740]};
ens0_layer0_N887 ens0_layer0_N887_inst (.M0(ens0_layer0_N887_wire), .M1(M1[887:887]));

wire [7:0] ens0_layer0_N888_wire = {M0[64], M0[80], M0[213], M0[291], M0[294], M0[571], M0[647], M0[712]};
ens0_layer0_N888 ens0_layer0_N888_inst (.M0(ens0_layer0_N888_wire), .M1(M1[888:888]));

wire [7:0] ens0_layer0_N889_wire = {M0[24], M0[144], M0[232], M0[355], M0[356], M0[386], M0[391], M0[570]};
ens0_layer0_N889 ens0_layer0_N889_inst (.M0(ens0_layer0_N889_wire), .M1(M1[889:889]));

wire [7:0] ens0_layer0_N890_wire = {M0[12], M0[162], M0[303], M0[325], M0[369], M0[630], M0[647], M0[761]};
ens0_layer0_N890 ens0_layer0_N890_inst (.M0(ens0_layer0_N890_wire), .M1(M1[890:890]));

wire [7:0] ens0_layer0_N891_wire = {M0[16], M0[19], M0[539], M0[569], M0[646], M0[701], M0[708], M0[714]};
ens0_layer0_N891 ens0_layer0_N891_inst (.M0(ens0_layer0_N891_wire), .M1(M1[891:891]));

wire [7:0] ens0_layer0_N892_wire = {M0[16], M0[23], M0[171], M0[214], M0[551], M0[576], M0[601], M0[774]};
ens0_layer0_N892 ens0_layer0_N892_inst (.M0(ens0_layer0_N892_wire), .M1(M1[892:892]));

wire [7:0] ens0_layer0_N893_wire = {M0[183], M0[311], M0[403], M0[413], M0[478], M0[524], M0[670], M0[721]};
ens0_layer0_N893 ens0_layer0_N893_inst (.M0(ens0_layer0_N893_wire), .M1(M1[893:893]));

wire [7:0] ens0_layer0_N894_wire = {M0[106], M0[216], M0[221], M0[482], M0[499], M0[692], M0[697], M0[723]};
ens0_layer0_N894 ens0_layer0_N894_inst (.M0(ens0_layer0_N894_wire), .M1(M1[894:894]));

wire [7:0] ens0_layer0_N895_wire = {M0[65], M0[129], M0[142], M0[163], M0[179], M0[182], M0[585], M0[706]};
ens0_layer0_N895 ens0_layer0_N895_inst (.M0(ens0_layer0_N895_wire), .M1(M1[895:895]));

wire [7:0] ens0_layer0_N896_wire = {M0[120], M0[448], M0[462], M0[554], M0[581], M0[593], M0[605], M0[629]};
ens0_layer0_N896 ens0_layer0_N896_inst (.M0(ens0_layer0_N896_wire), .M1(M1[896:896]));

wire [7:0] ens0_layer0_N897_wire = {M0[109], M0[232], M0[302], M0[404], M0[631], M0[685], M0[713], M0[775]};
ens0_layer0_N897 ens0_layer0_N897_inst (.M0(ens0_layer0_N897_wire), .M1(M1[897:897]));

wire [7:0] ens0_layer0_N898_wire = {M0[201], M0[205], M0[258], M0[274], M0[325], M0[483], M0[592], M0[607]};
ens0_layer0_N898 ens0_layer0_N898_inst (.M0(ens0_layer0_N898_wire), .M1(M1[898:898]));

wire [7:0] ens0_layer0_N899_wire = {M0[21], M0[67], M0[133], M0[184], M0[220], M0[462], M0[538], M0[603]};
ens0_layer0_N899 ens0_layer0_N899_inst (.M0(ens0_layer0_N899_wire), .M1(M1[899:899]));

wire [7:0] ens0_layer0_N900_wire = {M0[6], M0[343], M0[350], M0[377], M0[416], M0[442], M0[548], M0[586]};
ens0_layer0_N900 ens0_layer0_N900_inst (.M0(ens0_layer0_N900_wire), .M1(M1[900:900]));

wire [7:0] ens0_layer0_N901_wire = {M0[129], M0[214], M0[359], M0[371], M0[555], M0[684], M0[758], M0[782]};
ens0_layer0_N901 ens0_layer0_N901_inst (.M0(ens0_layer0_N901_wire), .M1(M1[901:901]));

wire [7:0] ens0_layer0_N902_wire = {M0[20], M0[195], M0[306], M0[384], M0[528], M0[608], M0[627], M0[638]};
ens0_layer0_N902 ens0_layer0_N902_inst (.M0(ens0_layer0_N902_wire), .M1(M1[902:902]));

wire [7:0] ens0_layer0_N903_wire = {M0[49], M0[392], M0[547], M0[576], M0[653], M0[680], M0[723], M0[772]};
ens0_layer0_N903 ens0_layer0_N903_inst (.M0(ens0_layer0_N903_wire), .M1(M1[903:903]));

wire [7:0] ens0_layer0_N904_wire = {M0[201], M0[253], M0[273], M0[347], M0[428], M0[442], M0[488], M0[592]};
ens0_layer0_N904 ens0_layer0_N904_inst (.M0(ens0_layer0_N904_wire), .M1(M1[904:904]));

wire [7:0] ens0_layer0_N905_wire = {M0[8], M0[258], M0[329], M0[340], M0[497], M0[619], M0[659], M0[727]};
ens0_layer0_N905 ens0_layer0_N905_inst (.M0(ens0_layer0_N905_wire), .M1(M1[905:905]));

wire [7:0] ens0_layer0_N906_wire = {M0[29], M0[88], M0[93], M0[123], M0[198], M0[552], M0[612], M0[670]};
ens0_layer0_N906 ens0_layer0_N906_inst (.M0(ens0_layer0_N906_wire), .M1(M1[906:906]));

wire [7:0] ens0_layer0_N907_wire = {M0[184], M0[294], M0[328], M0[338], M0[355], M0[515], M0[569], M0[694]};
ens0_layer0_N907 ens0_layer0_N907_inst (.M0(ens0_layer0_N907_wire), .M1(M1[907:907]));

wire [7:0] ens0_layer0_N908_wire = {M0[139], M0[332], M0[381], M0[388], M0[575], M0[595], M0[727], M0[766]};
ens0_layer0_N908 ens0_layer0_N908_inst (.M0(ens0_layer0_N908_wire), .M1(M1[908:908]));

wire [7:0] ens0_layer0_N909_wire = {M0[16], M0[113], M0[321], M0[367], M0[427], M0[677], M0[695], M0[697]};
ens0_layer0_N909 ens0_layer0_N909_inst (.M0(ens0_layer0_N909_wire), .M1(M1[909:909]));

wire [7:0] ens0_layer0_N910_wire = {M0[179], M0[404], M0[465], M0[490], M0[611], M0[619], M0[658], M0[767]};
ens0_layer0_N910 ens0_layer0_N910_inst (.M0(ens0_layer0_N910_wire), .M1(M1[910:910]));

wire [7:0] ens0_layer0_N911_wire = {M0[94], M0[255], M0[432], M0[546], M0[647], M0[669], M0[702], M0[768]};
ens0_layer0_N911 ens0_layer0_N911_inst (.M0(ens0_layer0_N911_wire), .M1(M1[911:911]));

wire [7:0] ens0_layer0_N912_wire = {M0[168], M0[198], M0[343], M0[446], M0[582], M0[687], M0[731], M0[783]};
ens0_layer0_N912 ens0_layer0_N912_inst (.M0(ens0_layer0_N912_wire), .M1(M1[912:912]));

wire [7:0] ens0_layer0_N913_wire = {M0[97], M0[216], M0[220], M0[490], M0[512], M0[545], M0[580], M0[783]};
ens0_layer0_N913 ens0_layer0_N913_inst (.M0(ens0_layer0_N913_wire), .M1(M1[913:913]));

wire [7:0] ens0_layer0_N914_wire = {M0[41], M0[55], M0[91], M0[116], M0[232], M0[380], M0[443], M0[637]};
ens0_layer0_N914 ens0_layer0_N914_inst (.M0(ens0_layer0_N914_wire), .M1(M1[914:914]));

wire [7:0] ens0_layer0_N915_wire = {M0[24], M0[81], M0[107], M0[199], M0[352], M0[427], M0[552], M0[782]};
ens0_layer0_N915 ens0_layer0_N915_inst (.M0(ens0_layer0_N915_wire), .M1(M1[915:915]));

wire [7:0] ens0_layer0_N916_wire = {M0[37], M0[92], M0[244], M0[293], M0[309], M0[424], M0[456], M0[562]};
ens0_layer0_N916 ens0_layer0_N916_inst (.M0(ens0_layer0_N916_wire), .M1(M1[916:916]));

wire [7:0] ens0_layer0_N917_wire = {M0[137], M0[155], M0[165], M0[539], M0[566], M0[634], M0[685], M0[781]};
ens0_layer0_N917 ens0_layer0_N917_inst (.M0(ens0_layer0_N917_wire), .M1(M1[917:917]));

wire [7:0] ens0_layer0_N918_wire = {M0[47], M0[147], M0[163], M0[257], M0[310], M0[315], M0[416], M0[540]};
ens0_layer0_N918 ens0_layer0_N918_inst (.M0(ens0_layer0_N918_wire), .M1(M1[918:918]));

wire [7:0] ens0_layer0_N919_wire = {M0[64], M0[245], M0[323], M0[369], M0[390], M0[532], M0[638], M0[686]};
ens0_layer0_N919 ens0_layer0_N919_inst (.M0(ens0_layer0_N919_wire), .M1(M1[919:919]));

wire [7:0] ens0_layer0_N920_wire = {M0[26], M0[132], M0[201], M0[426], M0[490], M0[546], M0[552], M0[747]};
ens0_layer0_N920 ens0_layer0_N920_inst (.M0(ens0_layer0_N920_wire), .M1(M1[920:920]));

wire [7:0] ens0_layer0_N921_wire = {M0[137], M0[269], M0[409], M0[432], M0[458], M0[538], M0[543], M0[742]};
ens0_layer0_N921 ens0_layer0_N921_inst (.M0(ens0_layer0_N921_wire), .M1(M1[921:921]));

wire [7:0] ens0_layer0_N922_wire = {M0[85], M0[197], M0[254], M0[321], M0[393], M0[634], M0[738], M0[775]};
ens0_layer0_N922 ens0_layer0_N922_inst (.M0(ens0_layer0_N922_wire), .M1(M1[922:922]));

wire [7:0] ens0_layer0_N923_wire = {M0[135], M0[286], M0[366], M0[426], M0[494], M0[672], M0[726], M0[761]};
ens0_layer0_N923 ens0_layer0_N923_inst (.M0(ens0_layer0_N923_wire), .M1(M1[923:923]));

wire [7:0] ens0_layer0_N924_wire = {M0[196], M0[249], M0[543], M0[547], M0[598], M0[602], M0[676], M0[680]};
ens0_layer0_N924 ens0_layer0_N924_inst (.M0(ens0_layer0_N924_wire), .M1(M1[924:924]));

wire [7:0] ens0_layer0_N925_wire = {M0[207], M0[331], M0[471], M0[600], M0[615], M0[616], M0[619], M0[766]};
ens0_layer0_N925 ens0_layer0_N925_inst (.M0(ens0_layer0_N925_wire), .M1(M1[925:925]));

wire [7:0] ens0_layer0_N926_wire = {M0[112], M0[289], M0[337], M0[433], M0[448], M0[520], M0[525], M0[724]};
ens0_layer0_N926 ens0_layer0_N926_inst (.M0(ens0_layer0_N926_wire), .M1(M1[926:926]));

wire [7:0] ens0_layer0_N927_wire = {M0[13], M0[223], M0[286], M0[318], M0[320], M0[603], M0[629], M0[747]};
ens0_layer0_N927 ens0_layer0_N927_inst (.M0(ens0_layer0_N927_wire), .M1(M1[927:927]));

wire [7:0] ens0_layer0_N928_wire = {M0[85], M0[102], M0[183], M0[215], M0[246], M0[292], M0[583], M0[636]};
ens0_layer0_N928 ens0_layer0_N928_inst (.M0(ens0_layer0_N928_wire), .M1(M1[928:928]));

wire [7:0] ens0_layer0_N929_wire = {M0[26], M0[164], M0[205], M0[223], M0[402], M0[528], M0[550], M0[686]};
ens0_layer0_N929 ens0_layer0_N929_inst (.M0(ens0_layer0_N929_wire), .M1(M1[929:929]));

wire [7:0] ens0_layer0_N930_wire = {M0[96], M0[294], M0[370], M0[437], M0[529], M0[530], M0[546], M0[712]};
ens0_layer0_N930 ens0_layer0_N930_inst (.M0(ens0_layer0_N930_wire), .M1(M1[930:930]));

wire [7:0] ens0_layer0_N931_wire = {M0[119], M0[159], M0[227], M0[347], M0[349], M0[369], M0[605], M0[769]};
ens0_layer0_N931 ens0_layer0_N931_inst (.M0(ens0_layer0_N931_wire), .M1(M1[931:931]));

wire [7:0] ens0_layer0_N932_wire = {M0[82], M0[117], M0[285], M0[287], M0[311], M0[417], M0[420], M0[570]};
ens0_layer0_N932 ens0_layer0_N932_inst (.M0(ens0_layer0_N932_wire), .M1(M1[932:932]));

wire [7:0] ens0_layer0_N933_wire = {M0[39], M0[194], M0[307], M0[368], M0[417], M0[422], M0[471], M0[557]};
ens0_layer0_N933 ens0_layer0_N933_inst (.M0(ens0_layer0_N933_wire), .M1(M1[933:933]));

wire [7:0] ens0_layer0_N934_wire = {M0[41], M0[145], M0[266], M0[460], M0[522], M0[556], M0[584], M0[778]};
ens0_layer0_N934 ens0_layer0_N934_inst (.M0(ens0_layer0_N934_wire), .M1(M1[934:934]));

wire [7:0] ens0_layer0_N935_wire = {M0[131], M0[399], M0[415], M0[464], M0[513], M0[515], M0[550], M0[597]};
ens0_layer0_N935 ens0_layer0_N935_inst (.M0(ens0_layer0_N935_wire), .M1(M1[935:935]));

wire [7:0] ens0_layer0_N936_wire = {M0[52], M0[138], M0[469], M0[534], M0[571], M0[700], M0[776], M0[780]};
ens0_layer0_N936 ens0_layer0_N936_inst (.M0(ens0_layer0_N936_wire), .M1(M1[936:936]));

wire [7:0] ens0_layer0_N937_wire = {M0[81], M0[191], M0[468], M0[549], M0[598], M0[611], M0[661], M0[694]};
ens0_layer0_N937 ens0_layer0_N937_inst (.M0(ens0_layer0_N937_wire), .M1(M1[937:937]));

wire [7:0] ens0_layer0_N938_wire = {M0[19], M0[121], M0[136], M0[175], M0[220], M0[370], M0[438], M0[523]};
ens0_layer0_N938 ens0_layer0_N938_inst (.M0(ens0_layer0_N938_wire), .M1(M1[938:938]));

wire [7:0] ens0_layer0_N939_wire = {M0[120], M0[185], M0[256], M0[359], M0[414], M0[491], M0[554], M0[762]};
ens0_layer0_N939 ens0_layer0_N939_inst (.M0(ens0_layer0_N939_wire), .M1(M1[939:939]));

wire [7:0] ens0_layer0_N940_wire = {M0[190], M0[369], M0[393], M0[436], M0[443], M0[444], M0[551], M0[556]};
ens0_layer0_N940 ens0_layer0_N940_inst (.M0(ens0_layer0_N940_wire), .M1(M1[940:940]));

wire [7:0] ens0_layer0_N941_wire = {M0[66], M0[445], M0[482], M0[594], M0[597], M0[656], M0[713], M0[783]};
ens0_layer0_N941 ens0_layer0_N941_inst (.M0(ens0_layer0_N941_wire), .M1(M1[941:941]));

wire [7:0] ens0_layer0_N942_wire = {M0[91], M0[297], M0[302], M0[342], M0[386], M0[409], M0[441], M0[749]};
ens0_layer0_N942 ens0_layer0_N942_inst (.M0(ens0_layer0_N942_wire), .M1(M1[942:942]));

wire [7:0] ens0_layer0_N943_wire = {M0[25], M0[95], M0[188], M0[288], M0[389], M0[444], M0[458], M0[482]};
ens0_layer0_N943 ens0_layer0_N943_inst (.M0(ens0_layer0_N943_wire), .M1(M1[943:943]));

wire [7:0] ens0_layer0_N944_wire = {M0[32], M0[190], M0[240], M0[256], M0[408], M0[529], M0[747], M0[751]};
ens0_layer0_N944 ens0_layer0_N944_inst (.M0(ens0_layer0_N944_wire), .M1(M1[944:944]));

wire [7:0] ens0_layer0_N945_wire = {M0[80], M0[209], M0[314], M0[332], M0[400], M0[436], M0[625], M0[705]};
ens0_layer0_N945 ens0_layer0_N945_inst (.M0(ens0_layer0_N945_wire), .M1(M1[945:945]));

wire [7:0] ens0_layer0_N946_wire = {M0[113], M0[277], M0[331], M0[390], M0[485], M0[563], M0[603], M0[719]};
ens0_layer0_N946 ens0_layer0_N946_inst (.M0(ens0_layer0_N946_wire), .M1(M1[946:946]));

wire [7:0] ens0_layer0_N947_wire = {M0[36], M0[133], M0[170], M0[206], M0[510], M0[557], M0[622], M0[746]};
ens0_layer0_N947 ens0_layer0_N947_inst (.M0(ens0_layer0_N947_wire), .M1(M1[947:947]));

wire [7:0] ens0_layer0_N948_wire = {M0[18], M0[157], M0[276], M0[492], M0[544], M0[580], M0[637], M0[737]};
ens0_layer0_N948 ens0_layer0_N948_inst (.M0(ens0_layer0_N948_wire), .M1(M1[948:948]));

wire [7:0] ens0_layer0_N949_wire = {M0[0], M0[54], M0[152], M0[163], M0[264], M0[284], M0[314], M0[525]};
ens0_layer0_N949 ens0_layer0_N949_inst (.M0(ens0_layer0_N949_wire), .M1(M1[949:949]));

wire [7:0] ens0_layer0_N950_wire = {M0[1], M0[43], M0[113], M0[307], M0[315], M0[448], M0[459], M0[699]};
ens0_layer0_N950 ens0_layer0_N950_inst (.M0(ens0_layer0_N950_wire), .M1(M1[950:950]));

wire [7:0] ens0_layer0_N951_wire = {M0[92], M0[237], M0[317], M0[501], M0[594], M0[690], M0[710], M0[776]};
ens0_layer0_N951 ens0_layer0_N951_inst (.M0(ens0_layer0_N951_wire), .M1(M1[951:951]));

wire [7:0] ens0_layer0_N952_wire = {M0[27], M0[70], M0[201], M0[238], M0[252], M0[373], M0[497], M0[677]};
ens0_layer0_N952 ens0_layer0_N952_inst (.M0(ens0_layer0_N952_wire), .M1(M1[952:952]));

wire [7:0] ens0_layer0_N953_wire = {M0[199], M0[200], M0[328], M0[438], M0[514], M0[529], M0[580], M0[610]};
ens0_layer0_N953 ens0_layer0_N953_inst (.M0(ens0_layer0_N953_wire), .M1(M1[953:953]));

wire [7:0] ens0_layer0_N954_wire = {M0[18], M0[292], M0[453], M0[533], M0[560], M0[571], M0[593], M0[782]};
ens0_layer0_N954 ens0_layer0_N954_inst (.M0(ens0_layer0_N954_wire), .M1(M1[954:954]));

wire [7:0] ens0_layer0_N955_wire = {M0[185], M0[193], M0[203], M0[406], M0[453], M0[572], M0[584], M0[762]};
ens0_layer0_N955 ens0_layer0_N955_inst (.M0(ens0_layer0_N955_wire), .M1(M1[955:955]));

wire [7:0] ens0_layer0_N956_wire = {M0[151], M0[221], M0[368], M0[447], M0[449], M0[677], M0[707], M0[744]};
ens0_layer0_N956 ens0_layer0_N956_inst (.M0(ens0_layer0_N956_wire), .M1(M1[956:956]));

wire [7:0] ens0_layer0_N957_wire = {M0[181], M0[401], M0[468], M0[542], M0[548], M0[560], M0[604], M0[666]};
ens0_layer0_N957 ens0_layer0_N957_inst (.M0(ens0_layer0_N957_wire), .M1(M1[957:957]));

wire [7:0] ens0_layer0_N958_wire = {M0[57], M0[92], M0[314], M0[453], M0[604], M0[618], M0[674], M0[777]};
ens0_layer0_N958 ens0_layer0_N958_inst (.M0(ens0_layer0_N958_wire), .M1(M1[958:958]));

wire [7:0] ens0_layer0_N959_wire = {M0[35], M0[59], M0[81], M0[189], M0[199], M0[346], M0[536], M0[579]};
ens0_layer0_N959 ens0_layer0_N959_inst (.M0(ens0_layer0_N959_wire), .M1(M1[959:959]));

wire [7:0] ens0_layer0_N960_wire = {M0[110], M0[117], M0[370], M0[606], M0[657], M0[675], M0[779], M0[781]};
ens0_layer0_N960 ens0_layer0_N960_inst (.M0(ens0_layer0_N960_wire), .M1(M1[960:960]));

wire [7:0] ens0_layer0_N961_wire = {M0[239], M0[319], M0[338], M0[531], M0[541], M0[616], M0[666], M0[773]};
ens0_layer0_N961 ens0_layer0_N961_inst (.M0(ens0_layer0_N961_wire), .M1(M1[961:961]));

wire [7:0] ens0_layer0_N962_wire = {M0[86], M0[94], M0[147], M0[155], M0[173], M0[436], M0[538], M0[775]};
ens0_layer0_N962 ens0_layer0_N962_inst (.M0(ens0_layer0_N962_wire), .M1(M1[962:962]));

wire [7:0] ens0_layer0_N963_wire = {M0[69], M0[127], M0[227], M0[282], M0[402], M0[476], M0[540], M0[648]};
ens0_layer0_N963 ens0_layer0_N963_inst (.M0(ens0_layer0_N963_wire), .M1(M1[963:963]));

wire [7:0] ens0_layer0_N964_wire = {M0[125], M0[171], M0[258], M0[303], M0[334], M0[392], M0[446], M0[452]};
ens0_layer0_N964 ens0_layer0_N964_inst (.M0(ens0_layer0_N964_wire), .M1(M1[964:964]));

wire [7:0] ens0_layer0_N965_wire = {M0[56], M0[164], M0[190], M0[336], M0[451], M0[457], M0[525], M0[690]};
ens0_layer0_N965 ens0_layer0_N965_inst (.M0(ens0_layer0_N965_wire), .M1(M1[965:965]));

wire [7:0] ens0_layer0_N966_wire = {M0[56], M0[402], M0[482], M0[496], M0[549], M0[550], M0[571], M0[644]};
ens0_layer0_N966 ens0_layer0_N966_inst (.M0(ens0_layer0_N966_wire), .M1(M1[966:966]));

wire [7:0] ens0_layer0_N967_wire = {M0[38], M0[90], M0[146], M0[325], M0[461], M0[578], M0[659], M0[724]};
ens0_layer0_N967 ens0_layer0_N967_inst (.M0(ens0_layer0_N967_wire), .M1(M1[967:967]));

wire [7:0] ens0_layer0_N968_wire = {M0[160], M0[179], M0[188], M0[480], M0[507], M0[645], M0[664], M0[691]};
ens0_layer0_N968 ens0_layer0_N968_inst (.M0(ens0_layer0_N968_wire), .M1(M1[968:968]));

wire [7:0] ens0_layer0_N969_wire = {M0[1], M0[44], M0[63], M0[99], M0[126], M0[312], M0[526], M0[704]};
ens0_layer0_N969 ens0_layer0_N969_inst (.M0(ens0_layer0_N969_wire), .M1(M1[969:969]));

wire [7:0] ens0_layer0_N970_wire = {M0[47], M0[56], M0[151], M0[203], M0[236], M0[249], M0[292], M0[383]};
ens0_layer0_N970 ens0_layer0_N970_inst (.M0(ens0_layer0_N970_wire), .M1(M1[970:970]));

wire [7:0] ens0_layer0_N971_wire = {M0[326], M0[431], M0[455], M0[494], M0[580], M0[590], M0[664], M0[735]};
ens0_layer0_N971 ens0_layer0_N971_inst (.M0(ens0_layer0_N971_wire), .M1(M1[971:971]));

wire [7:0] ens0_layer0_N972_wire = {M0[79], M0[130], M0[238], M0[336], M0[421], M0[440], M0[486], M0[593]};
ens0_layer0_N972 ens0_layer0_N972_inst (.M0(ens0_layer0_N972_wire), .M1(M1[972:972]));

wire [7:0] ens0_layer0_N973_wire = {M0[165], M0[171], M0[222], M0[396], M0[451], M0[691], M0[712], M0[722]};
ens0_layer0_N973 ens0_layer0_N973_inst (.M0(ens0_layer0_N973_wire), .M1(M1[973:973]));

wire [7:0] ens0_layer0_N974_wire = {M0[167], M0[609], M0[686], M0[708], M0[731], M0[766], M0[782], M0[783]};
ens0_layer0_N974 ens0_layer0_N974_inst (.M0(ens0_layer0_N974_wire), .M1(M1[974:974]));

wire [7:0] ens0_layer0_N975_wire = {M0[55], M0[120], M0[202], M0[318], M0[354], M0[551], M0[615], M0[724]};
ens0_layer0_N975 ens0_layer0_N975_inst (.M0(ens0_layer0_N975_wire), .M1(M1[975:975]));

wire [7:0] ens0_layer0_N976_wire = {M0[41], M0[235], M0[261], M0[546], M0[569], M0[689], M0[749], M0[766]};
ens0_layer0_N976 ens0_layer0_N976_inst (.M0(ens0_layer0_N976_wire), .M1(M1[976:976]));

wire [7:0] ens0_layer0_N977_wire = {M0[31], M0[157], M0[172], M0[216], M0[222], M0[377], M0[645], M0[688]};
ens0_layer0_N977 ens0_layer0_N977_inst (.M0(ens0_layer0_N977_wire), .M1(M1[977:977]));

wire [7:0] ens0_layer0_N978_wire = {M0[33], M0[115], M0[153], M0[538], M0[616], M0[632], M0[760], M0[762]};
ens0_layer0_N978 ens0_layer0_N978_inst (.M0(ens0_layer0_N978_wire), .M1(M1[978:978]));

wire [7:0] ens0_layer0_N979_wire = {M0[17], M0[36], M0[265], M0[386], M0[453], M0[534], M0[609], M0[781]};
ens0_layer0_N979 ens0_layer0_N979_inst (.M0(ens0_layer0_N979_wire), .M1(M1[979:979]));

wire [7:0] ens0_layer0_N980_wire = {M0[25], M0[256], M0[333], M0[498], M0[586], M0[597], M0[633], M0[750]};
ens0_layer0_N980 ens0_layer0_N980_inst (.M0(ens0_layer0_N980_wire), .M1(M1[980:980]));

wire [7:0] ens0_layer0_N981_wire = {M0[5], M0[9], M0[176], M0[231], M0[519], M0[542], M0[680], M0[728]};
ens0_layer0_N981 ens0_layer0_N981_inst (.M0(ens0_layer0_N981_wire), .M1(M1[981:981]));

wire [7:0] ens0_layer0_N982_wire = {M0[99], M0[139], M0[177], M0[422], M0[452], M0[574], M0[618], M0[781]};
ens0_layer0_N982 ens0_layer0_N982_inst (.M0(ens0_layer0_N982_wire), .M1(M1[982:982]));

wire [7:0] ens0_layer0_N983_wire = {M0[40], M0[68], M0[210], M0[270], M0[349], M0[419], M0[585], M0[702]};
ens0_layer0_N983 ens0_layer0_N983_inst (.M0(ens0_layer0_N983_wire), .M1(M1[983:983]));

wire [7:0] ens0_layer0_N984_wire = {M0[13], M0[208], M0[258], M0[366], M0[540], M0[567], M0[590], M0[662]};
ens0_layer0_N984 ens0_layer0_N984_inst (.M0(ens0_layer0_N984_wire), .M1(M1[984:984]));

wire [7:0] ens0_layer0_N985_wire = {M0[15], M0[126], M0[132], M0[219], M0[277], M0[596], M0[654], M0[748]};
ens0_layer0_N985 ens0_layer0_N985_inst (.M0(ens0_layer0_N985_wire), .M1(M1[985:985]));

wire [7:0] ens0_layer0_N986_wire = {M0[57], M0[143], M0[326], M0[346], M0[413], M0[606], M0[644], M0[739]};
ens0_layer0_N986 ens0_layer0_N986_inst (.M0(ens0_layer0_N986_wire), .M1(M1[986:986]));

wire [7:0] ens0_layer0_N987_wire = {M0[50], M0[179], M0[202], M0[249], M0[324], M0[533], M0[564], M0[764]};
ens0_layer0_N987 ens0_layer0_N987_inst (.M0(ens0_layer0_N987_wire), .M1(M1[987:987]));

wire [7:0] ens0_layer0_N988_wire = {M0[133], M0[226], M0[509], M0[510], M0[561], M0[612], M0[622], M0[765]};
ens0_layer0_N988 ens0_layer0_N988_inst (.M0(ens0_layer0_N988_wire), .M1(M1[988:988]));

wire [7:0] ens0_layer0_N989_wire = {M0[166], M0[210], M0[272], M0[314], M0[467], M0[505], M0[536], M0[568]};
ens0_layer0_N989 ens0_layer0_N989_inst (.M0(ens0_layer0_N989_wire), .M1(M1[989:989]));

wire [7:0] ens0_layer0_N990_wire = {M0[302], M0[444], M0[476], M0[492], M0[494], M0[569], M0[749], M0[755]};
ens0_layer0_N990 ens0_layer0_N990_inst (.M0(ens0_layer0_N990_wire), .M1(M1[990:990]));

wire [7:0] ens0_layer0_N991_wire = {M0[47], M0[94], M0[120], M0[327], M0[405], M0[411], M0[710], M0[720]};
ens0_layer0_N991 ens0_layer0_N991_inst (.M0(ens0_layer0_N991_wire), .M1(M1[991:991]));

wire [7:0] ens0_layer0_N992_wire = {M0[22], M0[309], M0[340], M0[376], M0[462], M0[534], M0[639], M0[662]};
ens0_layer0_N992 ens0_layer0_N992_inst (.M0(ens0_layer0_N992_wire), .M1(M1[992:992]));

wire [7:0] ens0_layer0_N993_wire = {M0[25], M0[66], M0[137], M0[251], M0[270], M0[284], M0[378], M0[475]};
ens0_layer0_N993 ens0_layer0_N993_inst (.M0(ens0_layer0_N993_wire), .M1(M1[993:993]));

wire [7:0] ens0_layer0_N994_wire = {M0[29], M0[73], M0[128], M0[188], M0[251], M0[315], M0[339], M0[390]};
ens0_layer0_N994 ens0_layer0_N994_inst (.M0(ens0_layer0_N994_wire), .M1(M1[994:994]));

wire [7:0] ens0_layer0_N995_wire = {M0[85], M0[96], M0[98], M0[131], M0[180], M0[190], M0[278], M0[771]};
ens0_layer0_N995 ens0_layer0_N995_inst (.M0(ens0_layer0_N995_wire), .M1(M1[995:995]));

wire [7:0] ens0_layer0_N996_wire = {M0[51], M0[77], M0[227], M0[414], M0[415], M0[422], M0[547], M0[735]};
ens0_layer0_N996 ens0_layer0_N996_inst (.M0(ens0_layer0_N996_wire), .M1(M1[996:996]));

wire [7:0] ens0_layer0_N997_wire = {M0[126], M0[253], M0[291], M0[331], M0[372], M0[554], M0[614], M0[726]};
ens0_layer0_N997 ens0_layer0_N997_inst (.M0(ens0_layer0_N997_wire), .M1(M1[997:997]));

wire [7:0] ens0_layer0_N998_wire = {M0[75], M0[310], M0[434], M0[484], M0[521], M0[527], M0[663], M0[689]};
ens0_layer0_N998 ens0_layer0_N998_inst (.M0(ens0_layer0_N998_wire), .M1(M1[998:998]));

wire [7:0] ens0_layer0_N999_wire = {M0[179], M0[377], M0[378], M0[499], M0[644], M0[723], M0[726], M0[767]};
ens0_layer0_N999 ens0_layer0_N999_inst (.M0(ens0_layer0_N999_wire), .M1(M1[999:999]));

wire [7:0] ens0_layer0_N1000_wire = {M0[105], M0[107], M0[146], M0[534], M0[561], M0[665], M0[676], M0[687]};
ens0_layer0_N1000 ens0_layer0_N1000_inst (.M0(ens0_layer0_N1000_wire), .M1(M1[1000:1000]));

wire [7:0] ens0_layer0_N1001_wire = {M0[97], M0[111], M0[239], M0[281], M0[326], M0[613], M0[715], M0[768]};
ens0_layer0_N1001 ens0_layer0_N1001_inst (.M0(ens0_layer0_N1001_wire), .M1(M1[1001:1001]));

wire [7:0] ens0_layer0_N1002_wire = {M0[132], M0[178], M0[305], M0[394], M0[599], M0[600], M0[630], M0[707]};
ens0_layer0_N1002 ens0_layer0_N1002_inst (.M0(ens0_layer0_N1002_wire), .M1(M1[1002:1002]));

wire [7:0] ens0_layer0_N1003_wire = {M0[222], M0[327], M0[335], M0[483], M0[490], M0[555], M0[584], M0[641]};
ens0_layer0_N1003 ens0_layer0_N1003_inst (.M0(ens0_layer0_N1003_wire), .M1(M1[1003:1003]));

wire [7:0] ens0_layer0_N1004_wire = {M0[242], M0[243], M0[309], M0[334], M0[482], M0[528], M0[661], M0[736]};
ens0_layer0_N1004 ens0_layer0_N1004_inst (.M0(ens0_layer0_N1004_wire), .M1(M1[1004:1004]));

wire [7:0] ens0_layer0_N1005_wire = {M0[46], M0[120], M0[303], M0[356], M0[407], M0[632], M0[708], M0[743]};
ens0_layer0_N1005 ens0_layer0_N1005_inst (.M0(ens0_layer0_N1005_wire), .M1(M1[1005:1005]));

wire [7:0] ens0_layer0_N1006_wire = {M0[33], M0[345], M0[482], M0[571], M0[586], M0[676], M0[730], M0[764]};
ens0_layer0_N1006 ens0_layer0_N1006_inst (.M0(ens0_layer0_N1006_wire), .M1(M1[1006:1006]));

wire [7:0] ens0_layer0_N1007_wire = {M0[281], M0[295], M0[440], M0[529], M0[538], M0[554], M0[650], M0[767]};
ens0_layer0_N1007 ens0_layer0_N1007_inst (.M0(ens0_layer0_N1007_wire), .M1(M1[1007:1007]));

wire [7:0] ens0_layer0_N1008_wire = {M0[175], M0[336], M0[362], M0[421], M0[516], M0[630], M0[770], M0[782]};
ens0_layer0_N1008 ens0_layer0_N1008_inst (.M0(ens0_layer0_N1008_wire), .M1(M1[1008:1008]));

wire [7:0] ens0_layer0_N1009_wire = {M0[68], M0[135], M0[293], M0[521], M0[564], M0[614], M0[631], M0[641]};
ens0_layer0_N1009 ens0_layer0_N1009_inst (.M0(ens0_layer0_N1009_wire), .M1(M1[1009:1009]));

wire [7:0] ens0_layer0_N1010_wire = {M0[12], M0[136], M0[333], M0[624], M0[626], M0[657], M0[665], M0[685]};
ens0_layer0_N1010 ens0_layer0_N1010_inst (.M0(ens0_layer0_N1010_wire), .M1(M1[1010:1010]));

wire [7:0] ens0_layer0_N1011_wire = {M0[116], M0[128], M0[310], M0[492], M0[597], M0[678], M0[696], M0[712]};
ens0_layer0_N1011 ens0_layer0_N1011_inst (.M0(ens0_layer0_N1011_wire), .M1(M1[1011:1011]));

wire [7:0] ens0_layer0_N1012_wire = {M0[80], M0[183], M0[257], M0[263], M0[315], M0[331], M0[554], M0[585]};
ens0_layer0_N1012 ens0_layer0_N1012_inst (.M0(ens0_layer0_N1012_wire), .M1(M1[1012:1012]));

wire [7:0] ens0_layer0_N1013_wire = {M0[171], M0[298], M0[327], M0[526], M0[536], M0[557], M0[567], M0[737]};
ens0_layer0_N1013 ens0_layer0_N1013_inst (.M0(ens0_layer0_N1013_wire), .M1(M1[1013:1013]));

wire [7:0] ens0_layer0_N1014_wire = {M0[162], M0[269], M0[328], M0[353], M0[364], M0[487], M0[663], M0[716]};
ens0_layer0_N1014 ens0_layer0_N1014_inst (.M0(ens0_layer0_N1014_wire), .M1(M1[1014:1014]));

wire [7:0] ens0_layer0_N1015_wire = {M0[95], M0[206], M0[210], M0[211], M0[251], M0[651], M0[734], M0[761]};
ens0_layer0_N1015 ens0_layer0_N1015_inst (.M0(ens0_layer0_N1015_wire), .M1(M1[1015:1015]));

wire [7:0] ens0_layer0_N1016_wire = {M0[33], M0[106], M0[107], M0[263], M0[287], M0[369], M0[419], M0[499]};
ens0_layer0_N1016 ens0_layer0_N1016_inst (.M0(ens0_layer0_N1016_wire), .M1(M1[1016:1016]));

wire [7:0] ens0_layer0_N1017_wire = {M0[50], M0[97], M0[164], M0[277], M0[309], M0[530], M0[584], M0[674]};
ens0_layer0_N1017 ens0_layer0_N1017_inst (.M0(ens0_layer0_N1017_wire), .M1(M1[1017:1017]));

wire [7:0] ens0_layer0_N1018_wire = {M0[67], M0[181], M0[261], M0[301], M0[361], M0[537], M0[626], M0[766]};
ens0_layer0_N1018 ens0_layer0_N1018_inst (.M0(ens0_layer0_N1018_wire), .M1(M1[1018:1018]));

wire [7:0] ens0_layer0_N1019_wire = {M0[26], M0[40], M0[102], M0[124], M0[204], M0[214], M0[299], M0[409]};
ens0_layer0_N1019 ens0_layer0_N1019_inst (.M0(ens0_layer0_N1019_wire), .M1(M1[1019:1019]));

wire [7:0] ens0_layer0_N1020_wire = {M0[103], M0[268], M0[368], M0[448], M0[570], M0[663], M0[718], M0[750]};
ens0_layer0_N1020 ens0_layer0_N1020_inst (.M0(ens0_layer0_N1020_wire), .M1(M1[1020:1020]));

wire [7:0] ens0_layer0_N1021_wire = {M0[165], M0[198], M0[296], M0[351], M0[517], M0[637], M0[649], M0[705]};
ens0_layer0_N1021 ens0_layer0_N1021_inst (.M0(ens0_layer0_N1021_wire), .M1(M1[1021:1021]));

wire [7:0] ens0_layer0_N1022_wire = {M0[62], M0[75], M0[137], M0[155], M0[170], M0[185], M0[328], M0[618]};
ens0_layer0_N1022 ens0_layer0_N1022_inst (.M0(ens0_layer0_N1022_wire), .M1(M1[1022:1022]));

wire [7:0] ens0_layer0_N1023_wire = {M0[19], M0[126], M0[146], M0[386], M0[388], M0[480], M0[577], M0[723]};
ens0_layer0_N1023 ens0_layer0_N1023_inst (.M0(ens0_layer0_N1023_wire), .M1(M1[1023:1023]));

endmodule