module ens0_layer5 (input [1023:0] M0, output [127:0] M1);

wire [7:0] ens0_layer5_N0_wire = {M0[326], M0[436], M0[662], M0[741], M0[748], M0[787], M0[878], M0[913]};
ens0_layer5_N0 ens0_layer5_N0_inst (.M0(ens0_layer5_N0_wire), .M1(M1[0:0]));

wire [7:0] ens0_layer5_N1_wire = {M0[100], M0[160], M0[178], M0[297], M0[365], M0[410], M0[447], M0[517]};
ens0_layer5_N1 ens0_layer5_N1_inst (.M0(ens0_layer5_N1_wire), .M1(M1[1:1]));

wire [7:0] ens0_layer5_N2_wire = {M0[0], M0[21], M0[338], M0[394], M0[413], M0[576], M0[754], M0[954]};
ens0_layer5_N2 ens0_layer5_N2_inst (.M0(ens0_layer5_N2_wire), .M1(M1[2:2]));

wire [7:0] ens0_layer5_N3_wire = {M0[160], M0[227], M0[583], M0[585], M0[641], M0[666], M0[752], M0[921]};
ens0_layer5_N3 ens0_layer5_N3_inst (.M0(ens0_layer5_N3_wire), .M1(M1[3:3]));

wire [7:0] ens0_layer5_N4_wire = {M0[21], M0[295], M0[590], M0[600], M0[838], M0[851], M0[865], M0[869]};
ens0_layer5_N4 ens0_layer5_N4_inst (.M0(ens0_layer5_N4_wire), .M1(M1[4:4]));

wire [7:0] ens0_layer5_N5_wire = {M0[38], M0[104], M0[205], M0[490], M0[548], M0[549], M0[551], M0[887]};
ens0_layer5_N5 ens0_layer5_N5_inst (.M0(ens0_layer5_N5_wire), .M1(M1[5:5]));

wire [7:0] ens0_layer5_N6_wire = {M0[43], M0[139], M0[250], M0[287], M0[453], M0[518], M0[522], M0[699]};
ens0_layer5_N6 ens0_layer5_N6_inst (.M0(ens0_layer5_N6_wire), .M1(M1[6:6]));

wire [7:0] ens0_layer5_N7_wire = {M0[110], M0[136], M0[159], M0[259], M0[382], M0[586], M0[687], M0[875]};
ens0_layer5_N7 ens0_layer5_N7_inst (.M0(ens0_layer5_N7_wire), .M1(M1[7:7]));

wire [7:0] ens0_layer5_N8_wire = {M0[88], M0[509], M0[607], M0[659], M0[778], M0[816], M0[912], M0[994]};
ens0_layer5_N8 ens0_layer5_N8_inst (.M0(ens0_layer5_N8_wire), .M1(M1[8:8]));

wire [7:0] ens0_layer5_N9_wire = {M0[160], M0[188], M0[451], M0[530], M0[672], M0[680], M0[691], M0[918]};
ens0_layer5_N9 ens0_layer5_N9_inst (.M0(ens0_layer5_N9_wire), .M1(M1[9:9]));

wire [7:0] ens0_layer5_N10_wire = {M0[350], M0[515], M0[570], M0[625], M0[642], M0[748], M0[757], M0[929]};
ens0_layer5_N10 ens0_layer5_N10_inst (.M0(ens0_layer5_N10_wire), .M1(M1[10:10]));

wire [7:0] ens0_layer5_N11_wire = {M0[62], M0[359], M0[389], M0[434], M0[724], M0[855], M0[907], M0[908]};
ens0_layer5_N11 ens0_layer5_N11_inst (.M0(ens0_layer5_N11_wire), .M1(M1[11:11]));

wire [7:0] ens0_layer5_N12_wire = {M0[227], M0[636], M0[669], M0[709], M0[763], M0[957], M0[1014], M0[1023]};
ens0_layer5_N12 ens0_layer5_N12_inst (.M0(ens0_layer5_N12_wire), .M1(M1[12:12]));

wire [7:0] ens0_layer5_N13_wire = {M0[197], M0[256], M0[280], M0[350], M0[543], M0[710], M0[815], M0[880]};
ens0_layer5_N13 ens0_layer5_N13_inst (.M0(ens0_layer5_N13_wire), .M1(M1[13:13]));

wire [7:0] ens0_layer5_N14_wire = {M0[266], M0[375], M0[539], M0[692], M0[818], M0[821], M0[963], M0[1023]};
ens0_layer5_N14 ens0_layer5_N14_inst (.M0(ens0_layer5_N14_wire), .M1(M1[14:14]));

wire [7:0] ens0_layer5_N15_wire = {M0[219], M0[484], M0[535], M0[553], M0[641], M0[742], M0[766], M0[904]};
ens0_layer5_N15 ens0_layer5_N15_inst (.M0(ens0_layer5_N15_wire), .M1(M1[15:15]));

wire [7:0] ens0_layer5_N16_wire = {M0[169], M0[178], M0[372], M0[642], M0[715], M0[885], M0[907], M0[975]};
ens0_layer5_N16 ens0_layer5_N16_inst (.M0(ens0_layer5_N16_wire), .M1(M1[16:16]));

wire [7:0] ens0_layer5_N17_wire = {M0[7], M0[24], M0[184], M0[236], M0[473], M0[519], M0[674], M0[788]};
ens0_layer5_N17 ens0_layer5_N17_inst (.M0(ens0_layer5_N17_wire), .M1(M1[17:17]));

wire [7:0] ens0_layer5_N18_wire = {M0[94], M0[144], M0[377], M0[429], M0[561], M0[597], M0[659], M0[771]};
ens0_layer5_N18 ens0_layer5_N18_inst (.M0(ens0_layer5_N18_wire), .M1(M1[18:18]));

wire [7:0] ens0_layer5_N19_wire = {M0[2], M0[88], M0[211], M0[467], M0[582], M0[786], M0[877], M0[892]};
ens0_layer5_N19 ens0_layer5_N19_inst (.M0(ens0_layer5_N19_wire), .M1(M1[19:19]));

wire [7:0] ens0_layer5_N20_wire = {M0[419], M0[480], M0[493], M0[688], M0[701], M0[776], M0[795], M0[887]};
ens0_layer5_N20 ens0_layer5_N20_inst (.M0(ens0_layer5_N20_wire), .M1(M1[20:20]));

wire [7:0] ens0_layer5_N21_wire = {M0[12], M0[216], M0[310], M0[524], M0[637], M0[952], M0[956], M0[1018]};
ens0_layer5_N21 ens0_layer5_N21_inst (.M0(ens0_layer5_N21_wire), .M1(M1[21:21]));

wire [7:0] ens0_layer5_N22_wire = {M0[67], M0[105], M0[310], M0[426], M0[681], M0[686], M0[834], M0[1004]};
ens0_layer5_N22 ens0_layer5_N22_inst (.M0(ens0_layer5_N22_wire), .M1(M1[22:22]));

wire [7:0] ens0_layer5_N23_wire = {M0[149], M0[222], M0[230], M0[299], M0[495], M0[818], M0[918], M0[940]};
ens0_layer5_N23 ens0_layer5_N23_inst (.M0(ens0_layer5_N23_wire), .M1(M1[23:23]));

wire [7:0] ens0_layer5_N24_wire = {M0[47], M0[103], M0[225], M0[252], M0[354], M0[493], M0[822], M0[853]};
ens0_layer5_N24 ens0_layer5_N24_inst (.M0(ens0_layer5_N24_wire), .M1(M1[24:24]));

wire [7:0] ens0_layer5_N25_wire = {M0[35], M0[243], M0[305], M0[635], M0[770], M0[870], M0[963], M0[1008]};
ens0_layer5_N25 ens0_layer5_N25_inst (.M0(ens0_layer5_N25_wire), .M1(M1[25:25]));

wire [7:0] ens0_layer5_N26_wire = {M0[78], M0[88], M0[145], M0[217], M0[385], M0[500], M0[546], M0[868]};
ens0_layer5_N26 ens0_layer5_N26_inst (.M0(ens0_layer5_N26_wire), .M1(M1[26:26]));

wire [7:0] ens0_layer5_N27_wire = {M0[4], M0[283], M0[378], M0[502], M0[514], M0[719], M0[799], M0[803]};
ens0_layer5_N27 ens0_layer5_N27_inst (.M0(ens0_layer5_N27_wire), .M1(M1[27:27]));

wire [7:0] ens0_layer5_N28_wire = {M0[30], M0[53], M0[370], M0[535], M0[575], M0[728], M0[831], M0[895]};
ens0_layer5_N28 ens0_layer5_N28_inst (.M0(ens0_layer5_N28_wire), .M1(M1[28:28]));

wire [7:0] ens0_layer5_N29_wire = {M0[49], M0[66], M0[103], M0[310], M0[361], M0[719], M0[846], M0[1007]};
ens0_layer5_N29 ens0_layer5_N29_inst (.M0(ens0_layer5_N29_wire), .M1(M1[29:29]));

wire [7:0] ens0_layer5_N30_wire = {M0[232], M0[343], M0[405], M0[594], M0[641], M0[657], M0[817], M0[1006]};
ens0_layer5_N30 ens0_layer5_N30_inst (.M0(ens0_layer5_N30_wire), .M1(M1[30:30]));

wire [7:0] ens0_layer5_N31_wire = {M0[47], M0[88], M0[212], M0[223], M0[332], M0[552], M0[717], M0[875]};
ens0_layer5_N31 ens0_layer5_N31_inst (.M0(ens0_layer5_N31_wire), .M1(M1[31:31]));

wire [7:0] ens0_layer5_N32_wire = {M0[13], M0[44], M0[306], M0[442], M0[493], M0[569], M0[866], M0[911]};
ens0_layer5_N32 ens0_layer5_N32_inst (.M0(ens0_layer5_N32_wire), .M1(M1[32:32]));

wire [7:0] ens0_layer5_N33_wire = {M0[234], M0[271], M0[343], M0[432], M0[555], M0[578], M0[595], M0[830]};
ens0_layer5_N33 ens0_layer5_N33_inst (.M0(ens0_layer5_N33_wire), .M1(M1[33:33]));

wire [7:0] ens0_layer5_N34_wire = {M0[265], M0[266], M0[438], M0[526], M0[617], M0[622], M0[669], M0[804]};
ens0_layer5_N34 ens0_layer5_N34_inst (.M0(ens0_layer5_N34_wire), .M1(M1[34:34]));

wire [7:0] ens0_layer5_N35_wire = {M0[0], M0[297], M0[493], M0[530], M0[568], M0[692], M0[880], M0[1013]};
ens0_layer5_N35 ens0_layer5_N35_inst (.M0(ens0_layer5_N35_wire), .M1(M1[35:35]));

wire [7:0] ens0_layer5_N36_wire = {M0[180], M0[304], M0[336], M0[377], M0[805], M0[892], M0[894], M0[982]};
ens0_layer5_N36 ens0_layer5_N36_inst (.M0(ens0_layer5_N36_wire), .M1(M1[36:36]));

wire [7:0] ens0_layer5_N37_wire = {M0[23], M0[181], M0[247], M0[579], M0[711], M0[905], M0[906], M0[947]};
ens0_layer5_N37 ens0_layer5_N37_inst (.M0(ens0_layer5_N37_wire), .M1(M1[37:37]));

wire [7:0] ens0_layer5_N38_wire = {M0[56], M0[65], M0[129], M0[159], M0[323], M0[365], M0[825], M0[846]};
ens0_layer5_N38 ens0_layer5_N38_inst (.M0(ens0_layer5_N38_wire), .M1(M1[38:38]));

wire [7:0] ens0_layer5_N39_wire = {M0[10], M0[273], M0[290], M0[454], M0[574], M0[757], M0[931], M0[964]};
ens0_layer5_N39 ens0_layer5_N39_inst (.M0(ens0_layer5_N39_wire), .M1(M1[39:39]));

wire [7:0] ens0_layer5_N40_wire = {M0[39], M0[148], M0[162], M0[576], M0[633], M0[774], M0[834], M0[1015]};
ens0_layer5_N40 ens0_layer5_N40_inst (.M0(ens0_layer5_N40_wire), .M1(M1[40:40]));

wire [7:0] ens0_layer5_N41_wire = {M0[44], M0[344], M0[379], M0[432], M0[493], M0[720], M0[911], M0[948]};
ens0_layer5_N41 ens0_layer5_N41_inst (.M0(ens0_layer5_N41_wire), .M1(M1[41:41]));

wire [7:0] ens0_layer5_N42_wire = {M0[74], M0[289], M0[310], M0[386], M0[587], M0[645], M0[812], M0[937]};
ens0_layer5_N42 ens0_layer5_N42_inst (.M0(ens0_layer5_N42_wire), .M1(M1[42:42]));

wire [7:0] ens0_layer5_N43_wire = {M0[106], M0[276], M0[501], M0[685], M0[699], M0[844], M0[849], M0[948]};
ens0_layer5_N43 ens0_layer5_N43_inst (.M0(ens0_layer5_N43_wire), .M1(M1[43:43]));

wire [7:0] ens0_layer5_N44_wire = {M0[7], M0[122], M0[339], M0[354], M0[361], M0[477], M0[516], M0[1021]};
ens0_layer5_N44 ens0_layer5_N44_inst (.M0(ens0_layer5_N44_wire), .M1(M1[44:44]));

wire [7:0] ens0_layer5_N45_wire = {M0[189], M0[193], M0[222], M0[370], M0[386], M0[424], M0[531], M0[941]};
ens0_layer5_N45 ens0_layer5_N45_inst (.M0(ens0_layer5_N45_wire), .M1(M1[45:45]));

wire [7:0] ens0_layer5_N46_wire = {M0[103], M0[213], M0[219], M0[226], M0[303], M0[459], M0[881], M0[991]};
ens0_layer5_N46 ens0_layer5_N46_inst (.M0(ens0_layer5_N46_wire), .M1(M1[46:46]));

wire [7:0] ens0_layer5_N47_wire = {M0[77], M0[81], M0[165], M0[368], M0[377], M0[611], M0[753], M0[777]};
ens0_layer5_N47 ens0_layer5_N47_inst (.M0(ens0_layer5_N47_wire), .M1(M1[47:47]));

wire [7:0] ens0_layer5_N48_wire = {M0[36], M0[93], M0[134], M0[266], M0[441], M0[783], M0[875], M0[1007]};
ens0_layer5_N48 ens0_layer5_N48_inst (.M0(ens0_layer5_N48_wire), .M1(M1[48:48]));

wire [7:0] ens0_layer5_N49_wire = {M0[311], M0[570], M0[593], M0[629], M0[804], M0[841], M0[944], M0[949]};
ens0_layer5_N49 ens0_layer5_N49_inst (.M0(ens0_layer5_N49_wire), .M1(M1[49:49]));

wire [7:0] ens0_layer5_N50_wire = {M0[34], M0[47], M0[85], M0[154], M0[214], M0[294], M0[567], M0[943]};
ens0_layer5_N50 ens0_layer5_N50_inst (.M0(ens0_layer5_N50_wire), .M1(M1[50:50]));

wire [7:0] ens0_layer5_N51_wire = {M0[161], M0[283], M0[390], M0[481], M0[581], M0[661], M0[844], M0[965]};
ens0_layer5_N51 ens0_layer5_N51_inst (.M0(ens0_layer5_N51_wire), .M1(M1[51:51]));

wire [7:0] ens0_layer5_N52_wire = {M0[9], M0[28], M0[125], M0[349], M0[567], M0[642], M0[727], M0[881]};
ens0_layer5_N52 ens0_layer5_N52_inst (.M0(ens0_layer5_N52_wire), .M1(M1[52:52]));

wire [7:0] ens0_layer5_N53_wire = {M0[240], M0[273], M0[334], M0[355], M0[484], M0[755], M0[766], M0[917]};
ens0_layer5_N53 ens0_layer5_N53_inst (.M0(ens0_layer5_N53_wire), .M1(M1[53:53]));

wire [7:0] ens0_layer5_N54_wire = {M0[223], M0[342], M0[399], M0[544], M0[796], M0[859], M0[908], M0[911]};
ens0_layer5_N54 ens0_layer5_N54_inst (.M0(ens0_layer5_N54_wire), .M1(M1[54:54]));

wire [7:0] ens0_layer5_N55_wire = {M0[43], M0[51], M0[124], M0[233], M0[350], M0[472], M0[961], M0[1010]};
ens0_layer5_N55 ens0_layer5_N55_inst (.M0(ens0_layer5_N55_wire), .M1(M1[55:55]));

wire [7:0] ens0_layer5_N56_wire = {M0[4], M0[35], M0[64], M0[252], M0[343], M0[652], M0[653], M0[1009]};
ens0_layer5_N56 ens0_layer5_N56_inst (.M0(ens0_layer5_N56_wire), .M1(M1[56:56]));

wire [7:0] ens0_layer5_N57_wire = {M0[310], M0[367], M0[370], M0[488], M0[492], M0[532], M0[538], M0[647]};
ens0_layer5_N57 ens0_layer5_N57_inst (.M0(ens0_layer5_N57_wire), .M1(M1[57:57]));

wire [7:0] ens0_layer5_N58_wire = {M0[102], M0[151], M0[181], M0[219], M0[320], M0[596], M0[634], M0[888]};
ens0_layer5_N58 ens0_layer5_N58_inst (.M0(ens0_layer5_N58_wire), .M1(M1[58:58]));

wire [7:0] ens0_layer5_N59_wire = {M0[59], M0[373], M0[423], M0[665], M0[760], M0[882], M0[921], M0[924]};
ens0_layer5_N59 ens0_layer5_N59_inst (.M0(ens0_layer5_N59_wire), .M1(M1[59:59]));

wire [7:0] ens0_layer5_N60_wire = {M0[67], M0[190], M0[216], M0[262], M0[265], M0[299], M0[424], M0[811]};
ens0_layer5_N60 ens0_layer5_N60_inst (.M0(ens0_layer5_N60_wire), .M1(M1[60:60]));

wire [7:0] ens0_layer5_N61_wire = {M0[204], M0[390], M0[542], M0[571], M0[596], M0[677], M0[796], M0[808]};
ens0_layer5_N61 ens0_layer5_N61_inst (.M0(ens0_layer5_N61_wire), .M1(M1[61:61]));

wire [7:0] ens0_layer5_N62_wire = {M0[136], M0[188], M0[201], M0[317], M0[526], M0[660], M0[685], M0[826]};
ens0_layer5_N62 ens0_layer5_N62_inst (.M0(ens0_layer5_N62_wire), .M1(M1[62:62]));

wire [7:0] ens0_layer5_N63_wire = {M0[130], M0[193], M0[514], M0[604], M0[607], M0[767], M0[868], M0[1020]};
ens0_layer5_N63 ens0_layer5_N63_inst (.M0(ens0_layer5_N63_wire), .M1(M1[63:63]));

wire [7:0] ens0_layer5_N64_wire = {M0[32], M0[327], M0[520], M0[630], M0[720], M0[725], M0[823], M0[942]};
ens0_layer5_N64 ens0_layer5_N64_inst (.M0(ens0_layer5_N64_wire), .M1(M1[64:64]));

wire [7:0] ens0_layer5_N65_wire = {M0[34], M0[215], M0[341], M0[461], M0[517], M0[521], M0[754], M0[898]};
ens0_layer5_N65 ens0_layer5_N65_inst (.M0(ens0_layer5_N65_wire), .M1(M1[65:65]));

wire [7:0] ens0_layer5_N66_wire = {M0[39], M0[63], M0[96], M0[110], M0[302], M0[395], M0[625], M0[802]};
ens0_layer5_N66 ens0_layer5_N66_inst (.M0(ens0_layer5_N66_wire), .M1(M1[66:66]));

wire [7:0] ens0_layer5_N67_wire = {M0[89], M0[217], M0[255], M0[374], M0[597], M0[668], M0[773], M0[958]};
ens0_layer5_N67 ens0_layer5_N67_inst (.M0(ens0_layer5_N67_wire), .M1(M1[67:67]));

wire [7:0] ens0_layer5_N68_wire = {M0[468], M0[542], M0[569], M0[775], M0[848], M0[855], M0[893], M0[918]};
ens0_layer5_N68 ens0_layer5_N68_inst (.M0(ens0_layer5_N68_wire), .M1(M1[68:68]));

wire [7:0] ens0_layer5_N69_wire = {M0[34], M0[122], M0[368], M0[500], M0[527], M0[694], M0[726], M0[862]};
ens0_layer5_N69 ens0_layer5_N69_inst (.M0(ens0_layer5_N69_wire), .M1(M1[69:69]));

wire [7:0] ens0_layer5_N70_wire = {M0[30], M0[151], M0[236], M0[524], M0[525], M0[738], M0[995], M0[1012]};
ens0_layer5_N70 ens0_layer5_N70_inst (.M0(ens0_layer5_N70_wire), .M1(M1[70:70]));

wire [7:0] ens0_layer5_N71_wire = {M0[73], M0[95], M0[129], M0[178], M0[365], M0[374], M0[569], M0[725]};
ens0_layer5_N71 ens0_layer5_N71_inst (.M0(ens0_layer5_N71_wire), .M1(M1[71:71]));

wire [7:0] ens0_layer5_N72_wire = {M0[199], M0[260], M0[293], M0[423], M0[529], M0[543], M0[893], M0[930]};
ens0_layer5_N72 ens0_layer5_N72_inst (.M0(ens0_layer5_N72_wire), .M1(M1[72:72]));

wire [7:0] ens0_layer5_N73_wire = {M0[112], M0[262], M0[303], M0[566], M0[657], M0[850], M0[918], M0[958]};
ens0_layer5_N73 ens0_layer5_N73_inst (.M0(ens0_layer5_N73_wire), .M1(M1[73:73]));

wire [7:0] ens0_layer5_N74_wire = {M0[65], M0[176], M0[208], M0[258], M0[458], M0[588], M0[806], M0[889]};
ens0_layer5_N74 ens0_layer5_N74_inst (.M0(ens0_layer5_N74_wire), .M1(M1[74:74]));

wire [7:0] ens0_layer5_N75_wire = {M0[54], M0[158], M0[269], M0[512], M0[700], M0[813], M0[968], M0[992]};
ens0_layer5_N75 ens0_layer5_N75_inst (.M0(ens0_layer5_N75_wire), .M1(M1[75:75]));

wire [7:0] ens0_layer5_N76_wire = {M0[78], M0[172], M0[319], M0[335], M0[514], M0[727], M0[736], M0[793]};
ens0_layer5_N76 ens0_layer5_N76_inst (.M0(ens0_layer5_N76_wire), .M1(M1[76:76]));

wire [7:0] ens0_layer5_N77_wire = {M0[92], M0[227], M0[254], M0[537], M0[585], M0[750], M0[914], M0[977]};
ens0_layer5_N77 ens0_layer5_N77_inst (.M0(ens0_layer5_N77_wire), .M1(M1[77:77]));

wire [7:0] ens0_layer5_N78_wire = {M0[224], M0[235], M0[286], M0[518], M0[702], M0[808], M0[840], M0[956]};
ens0_layer5_N78 ens0_layer5_N78_inst (.M0(ens0_layer5_N78_wire), .M1(M1[78:78]));

wire [7:0] ens0_layer5_N79_wire = {M0[99], M0[128], M0[142], M0[294], M0[376], M0[750], M0[899], M0[979]};
ens0_layer5_N79 ens0_layer5_N79_inst (.M0(ens0_layer5_N79_wire), .M1(M1[79:79]));

wire [7:0] ens0_layer5_N80_wire = {M0[118], M0[141], M0[385], M0[386], M0[501], M0[730], M0[789], M0[829]};
ens0_layer5_N80 ens0_layer5_N80_inst (.M0(ens0_layer5_N80_wire), .M1(M1[80:80]));

wire [7:0] ens0_layer5_N81_wire = {M0[169], M0[208], M0[258], M0[426], M0[611], M0[686], M0[876], M0[894]};
ens0_layer5_N81 ens0_layer5_N81_inst (.M0(ens0_layer5_N81_wire), .M1(M1[81:81]));

wire [7:0] ens0_layer5_N82_wire = {M0[175], M0[276], M0[464], M0[539], M0[558], M0[560], M0[567], M0[704]};
ens0_layer5_N82 ens0_layer5_N82_inst (.M0(ens0_layer5_N82_wire), .M1(M1[82:82]));

wire [7:0] ens0_layer5_N83_wire = {M0[90], M0[236], M0[250], M0[791], M0[834], M0[855], M0[967], M0[999]};
ens0_layer5_N83 ens0_layer5_N83_inst (.M0(ens0_layer5_N83_wire), .M1(M1[83:83]));

wire [7:0] ens0_layer5_N84_wire = {M0[101], M0[259], M0[267], M0[303], M0[632], M0[642], M0[872], M0[954]};
ens0_layer5_N84 ens0_layer5_N84_inst (.M0(ens0_layer5_N84_wire), .M1(M1[84:84]));

wire [7:0] ens0_layer5_N85_wire = {M0[97], M0[311], M0[430], M0[637], M0[706], M0[720], M0[738], M0[739]};
ens0_layer5_N85 ens0_layer5_N85_inst (.M0(ens0_layer5_N85_wire), .M1(M1[85:85]));

wire [7:0] ens0_layer5_N86_wire = {M0[172], M0[352], M0[460], M0[637], M0[814], M0[815], M0[905], M0[989]};
ens0_layer5_N86 ens0_layer5_N86_inst (.M0(ens0_layer5_N86_wire), .M1(M1[86:86]));

wire [7:0] ens0_layer5_N87_wire = {M0[52], M0[62], M0[306], M0[574], M0[589], M0[667], M0[828], M0[986]};
ens0_layer5_N87 ens0_layer5_N87_inst (.M0(ens0_layer5_N87_wire), .M1(M1[87:87]));

wire [7:0] ens0_layer5_N88_wire = {M0[6], M0[40], M0[187], M0[390], M0[738], M0[888], M0[957], M0[1022]};
ens0_layer5_N88 ens0_layer5_N88_inst (.M0(ens0_layer5_N88_wire), .M1(M1[88:88]));

wire [7:0] ens0_layer5_N89_wire = {M0[25], M0[63], M0[436], M0[537], M0[555], M0[597], M0[988], M0[1010]};
ens0_layer5_N89 ens0_layer5_N89_inst (.M0(ens0_layer5_N89_wire), .M1(M1[89:89]));

wire [7:0] ens0_layer5_N90_wire = {M0[221], M0[253], M0[304], M0[505], M0[581], M0[680], M0[699], M0[982]};
ens0_layer5_N90 ens0_layer5_N90_inst (.M0(ens0_layer5_N90_wire), .M1(M1[90:90]));

wire [7:0] ens0_layer5_N91_wire = {M0[3], M0[405], M0[441], M0[475], M0[530], M0[535], M0[748], M0[967]};
ens0_layer5_N91 ens0_layer5_N91_inst (.M0(ens0_layer5_N91_wire), .M1(M1[91:91]));

wire [7:0] ens0_layer5_N92_wire = {M0[67], M0[252], M0[378], M0[450], M0[510], M0[772], M0[806], M0[874]};
ens0_layer5_N92 ens0_layer5_N92_inst (.M0(ens0_layer5_N92_wire), .M1(M1[92:92]));

wire [7:0] ens0_layer5_N93_wire = {M0[16], M0[140], M0[211], M0[336], M0[465], M0[677], M0[746], M0[934]};
ens0_layer5_N93 ens0_layer5_N93_inst (.M0(ens0_layer5_N93_wire), .M1(M1[93:93]));

wire [7:0] ens0_layer5_N94_wire = {M0[5], M0[7], M0[135], M0[333], M0[380], M0[395], M0[610], M0[712]};
ens0_layer5_N94 ens0_layer5_N94_inst (.M0(ens0_layer5_N94_wire), .M1(M1[94:94]));

wire [7:0] ens0_layer5_N95_wire = {M0[249], M0[385], M0[407], M0[485], M0[602], M0[639], M0[816], M0[854]};
ens0_layer5_N95 ens0_layer5_N95_inst (.M0(ens0_layer5_N95_wire), .M1(M1[95:95]));

wire [7:0] ens0_layer5_N96_wire = {M0[60], M0[75], M0[424], M0[469], M0[694], M0[749], M0[792], M0[892]};
ens0_layer5_N96 ens0_layer5_N96_inst (.M0(ens0_layer5_N96_wire), .M1(M1[96:96]));

wire [7:0] ens0_layer5_N97_wire = {M0[347], M0[399], M0[689], M0[738], M0[846], M0[925], M0[941], M0[956]};
ens0_layer5_N97 ens0_layer5_N97_inst (.M0(ens0_layer5_N97_wire), .M1(M1[97:97]));

wire [7:0] ens0_layer5_N98_wire = {M0[81], M0[428], M0[467], M0[488], M0[640], M0[664], M0[862], M0[970]};
ens0_layer5_N98 ens0_layer5_N98_inst (.M0(ens0_layer5_N98_wire), .M1(M1[98:98]));

wire [7:0] ens0_layer5_N99_wire = {M0[97], M0[120], M0[195], M0[265], M0[603], M0[757], M0[870], M0[901]};
ens0_layer5_N99 ens0_layer5_N99_inst (.M0(ens0_layer5_N99_wire), .M1(M1[99:99]));

wire [7:0] ens0_layer5_N100_wire = {M0[118], M0[236], M0[393], M0[485], M0[543], M0[775], M0[820], M0[858]};
ens0_layer5_N100 ens0_layer5_N100_inst (.M0(ens0_layer5_N100_wire), .M1(M1[100:100]));

wire [7:0] ens0_layer5_N101_wire = {M0[7], M0[207], M0[208], M0[263], M0[268], M0[412], M0[490], M0[614]};
ens0_layer5_N101 ens0_layer5_N101_inst (.M0(ens0_layer5_N101_wire), .M1(M1[101:101]));

wire [7:0] ens0_layer5_N102_wire = {M0[6], M0[350], M0[354], M0[515], M0[622], M0[879], M0[914], M0[963]};
ens0_layer5_N102 ens0_layer5_N102_inst (.M0(ens0_layer5_N102_wire), .M1(M1[102:102]));

wire [7:0] ens0_layer5_N103_wire = {M0[49], M0[238], M0[374], M0[536], M0[613], M0[617], M0[791], M0[807]};
ens0_layer5_N103 ens0_layer5_N103_inst (.M0(ens0_layer5_N103_wire), .M1(M1[103:103]));

wire [7:0] ens0_layer5_N104_wire = {M0[139], M0[318], M0[405], M0[507], M0[621], M0[672], M0[818], M0[973]};
ens0_layer5_N104 ens0_layer5_N104_inst (.M0(ens0_layer5_N104_wire), .M1(M1[104:104]));

wire [7:0] ens0_layer5_N105_wire = {M0[72], M0[113], M0[168], M0[294], M0[436], M0[679], M0[700], M0[996]};
ens0_layer5_N105 ens0_layer5_N105_inst (.M0(ens0_layer5_N105_wire), .M1(M1[105:105]));

wire [7:0] ens0_layer5_N106_wire = {M0[300], M0[311], M0[441], M0[445], M0[678], M0[714], M0[905], M0[999]};
ens0_layer5_N106 ens0_layer5_N106_inst (.M0(ens0_layer5_N106_wire), .M1(M1[106:106]));

wire [7:0] ens0_layer5_N107_wire = {M0[59], M0[201], M0[456], M0[461], M0[522], M0[670], M0[732], M0[984]};
ens0_layer5_N107 ens0_layer5_N107_inst (.M0(ens0_layer5_N107_wire), .M1(M1[107:107]));

wire [7:0] ens0_layer5_N108_wire = {M0[402], M0[448], M0[452], M0[676], M0[789], M0[798], M0[834], M0[853]};
ens0_layer5_N108 ens0_layer5_N108_inst (.M0(ens0_layer5_N108_wire), .M1(M1[108:108]));

wire [7:0] ens0_layer5_N109_wire = {M0[125], M0[159], M0[221], M0[315], M0[378], M0[657], M0[777], M0[823]};
ens0_layer5_N109 ens0_layer5_N109_inst (.M0(ens0_layer5_N109_wire), .M1(M1[109:109]));

wire [7:0] ens0_layer5_N110_wire = {M0[40], M0[181], M0[203], M0[399], M0[439], M0[671], M0[897], M0[916]};
ens0_layer5_N110 ens0_layer5_N110_inst (.M0(ens0_layer5_N110_wire), .M1(M1[110:110]));

wire [7:0] ens0_layer5_N111_wire = {M0[144], M0[172], M0[364], M0[451], M0[604], M0[655], M0[874], M0[947]};
ens0_layer5_N111 ens0_layer5_N111_inst (.M0(ens0_layer5_N111_wire), .M1(M1[111:111]));

wire [7:0] ens0_layer5_N112_wire = {M0[71], M0[163], M0[197], M0[265], M0[331], M0[430], M0[852], M0[879]};
ens0_layer5_N112 ens0_layer5_N112_inst (.M0(ens0_layer5_N112_wire), .M1(M1[112:112]));

wire [7:0] ens0_layer5_N113_wire = {M0[69], M0[221], M0[463], M0[670], M0[680], M0[791], M0[811], M0[876]};
ens0_layer5_N113 ens0_layer5_N113_inst (.M0(ens0_layer5_N113_wire), .M1(M1[113:113]));

wire [7:0] ens0_layer5_N114_wire = {M0[24], M0[144], M0[283], M0[349], M0[389], M0[470], M0[508], M0[851]};
ens0_layer5_N114 ens0_layer5_N114_inst (.M0(ens0_layer5_N114_wire), .M1(M1[114:114]));

wire [7:0] ens0_layer5_N115_wire = {M0[131], M0[169], M0[210], M0[420], M0[537], M0[545], M0[618], M0[853]};
ens0_layer5_N115 ens0_layer5_N115_inst (.M0(ens0_layer5_N115_wire), .M1(M1[115:115]));

wire [7:0] ens0_layer5_N116_wire = {M0[446], M0[453], M0[517], M0[556], M0[868], M0[944], M0[958], M0[1010]};
ens0_layer5_N116 ens0_layer5_N116_inst (.M0(ens0_layer5_N116_wire), .M1(M1[116:116]));

wire [7:0] ens0_layer5_N117_wire = {M0[237], M0[344], M0[415], M0[486], M0[612], M0[847], M0[856], M0[941]};
ens0_layer5_N117 ens0_layer5_N117_inst (.M0(ens0_layer5_N117_wire), .M1(M1[117:117]));

wire [7:0] ens0_layer5_N118_wire = {M0[58], M0[317], M0[406], M0[460], M0[588], M0[697], M0[757], M0[1006]};
ens0_layer5_N118 ens0_layer5_N118_inst (.M0(ens0_layer5_N118_wire), .M1(M1[118:118]));

wire [7:0] ens0_layer5_N119_wire = {M0[151], M0[326], M0[459], M0[698], M0[704], M0[827], M0[927], M0[985]};
ens0_layer5_N119 ens0_layer5_N119_inst (.M0(ens0_layer5_N119_wire), .M1(M1[119:119]));

wire [7:0] ens0_layer5_N120_wire = {M0[12], M0[155], M0[275], M0[281], M0[433], M0[648], M0[802], M0[832]};
ens0_layer5_N120 ens0_layer5_N120_inst (.M0(ens0_layer5_N120_wire), .M1(M1[120:120]));

wire [7:0] ens0_layer5_N121_wire = {M0[23], M0[79], M0[165], M0[214], M0[362], M0[819], M0[943], M0[965]};
ens0_layer5_N121 ens0_layer5_N121_inst (.M0(ens0_layer5_N121_wire), .M1(M1[121:121]));

wire [7:0] ens0_layer5_N122_wire = {M0[140], M0[171], M0[317], M0[361], M0[371], M0[653], M0[773], M0[1001]};
ens0_layer5_N122 ens0_layer5_N122_inst (.M0(ens0_layer5_N122_wire), .M1(M1[122:122]));

wire [7:0] ens0_layer5_N123_wire = {M0[83], M0[95], M0[181], M0[207], M0[690], M0[819], M0[842], M0[913]};
ens0_layer5_N123 ens0_layer5_N123_inst (.M0(ens0_layer5_N123_wire), .M1(M1[123:123]));

wire [7:0] ens0_layer5_N124_wire = {M0[45], M0[203], M0[225], M0[387], M0[425], M0[767], M0[801], M0[916]};
ens0_layer5_N124 ens0_layer5_N124_inst (.M0(ens0_layer5_N124_wire), .M1(M1[124:124]));

wire [7:0] ens0_layer5_N125_wire = {M0[142], M0[189], M0[296], M0[451], M0[536], M0[810], M0[936], M0[952]};
ens0_layer5_N125 ens0_layer5_N125_inst (.M0(ens0_layer5_N125_wire), .M1(M1[125:125]));

wire [7:0] ens0_layer5_N126_wire = {M0[113], M0[253], M0[259], M0[304], M0[427], M0[644], M0[934], M0[974]};
ens0_layer5_N126 ens0_layer5_N126_inst (.M0(ens0_layer5_N126_wire), .M1(M1[126:126]));

wire [7:0] ens0_layer5_N127_wire = {M0[158], M0[208], M0[247], M0[632], M0[633], M0[661], M0[752], M0[958]};
ens0_layer5_N127 ens0_layer5_N127_inst (.M0(ens0_layer5_N127_wire), .M1(M1[127:127]));

endmodule